��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� j^ꘜI��e�cA�l�eף@�M����s�v��7-�1����P{A�2������J�ݮ�F�!ԪdX>��$aL�nHFig([䩾�Wj0�g��@i�*�E�ع�������x�f�Κ)���9]C��p�p���M7\����}m�����B��H��2�Md��])\ΤV\:�n5R�#Ӈ����,sdymK���������`*e;�Lɡ8�;��P��[�iΝ)Z�gQ�ƉJM]>��ő(�[�wO����X�,6L��f�Py�Jo"��aɗ栴�� ���x�5G�1?A����iǫa]r�YH���uh>� �W ��}�W��LI�j����\SQE��u�U^N�bbW]ަ���� R�8��FrO~jB��h�q�/'�51��-/�ϳz�B��=p-�������Zax����ʙ[N��1���(j,���W8�[b��V�:��-�L��5����zaF����ʿty�����I,^n#p)ˉZ��U�P7�AD��J�>&���mư='1O~����{��` ��v����a9D��c�gm����H~f�����a�=��P��!.od4|G�I��Cg̤y��@��۞/%�����h�c��5K�����{;K��AC�x�ӱX�"p�nXQ�&�n ��D2G=]�x��3�����=?���H̯R<QK����(����GZy^s������Y���y��%�ed�jKhXwxǮ�RKX��}���ι2r�Ãv�ĳG<ށ�sl�s8B�4� ��Qz2`�6��7����C��g�}�6>���n\:�^O�Vsz9T�׋u���� A�2(�q�+�H��#8�d���J� �ߜ87��kj$���!��ߩ(�«g�.�(0���f�[F�e�{��ey�`�C���A�d�7�!���7A�G��{�����:�{�M�d���X����<X�*D!���s�LGJ!��ba�.���L�r5�cKN���DGAm����K�k&j?%'��k�t2@+���*�M�vٔ ?6����V�C��h{�2�	y��`OF4#5wZl�͏E%�|�7 :f������Y��=�.Mpk|Tth w�c�`��c���+b��3~hqD�~!5��V���������~}���@��Ů���Ѣ�eJzϧhbGr(ȱ�����x�L�g.��Dc�R,� K9��/�	���F{�ꞷ%=�  �0|�H�ъ�n�ٗc�0hO/���~t�۬%�����U�`���)zR��>�=�;>n����d��c��#S��b���I�9��:33䄆��R
�S���꜇�2]��.KL%��U{AΉ�V�W��@5+��r������H&m ����0T|4��p�*Q�d�����*LO:�|k�W��5��t<��Mn�z`xǵ�Ɨ%
�q́�����UL�;2G���zS��9�x��Fa�~��31I�:�c剝���H$-vӑ�{l�{v �O�N:�P�{�`���,w�q��L�Ho�`�gFk��A�n�:�B�F5���	V1���'� %���������������WG�J�Lp؁5��Õ����N�I��+F���7	���}�*(BT��|"�W퀯[|"�J�s�D��?��{�%W0�}��m#�KU��bO��Rv�(C �ʾTfTiL�L��hDlD��G�+I���Z�RW V�(�7F2-h���!����z�P]j���]}��v�Z���n��Xǁ`3B�Z�vN{b M �t*��͆s�̳�R�_?��$�P���&SN�]p�]蒦���w���ƨ�̵z�9��K��,\�h�%x��$Q�a7Jr���x�K1 ��k�*�����(���QةLx�tît�3�ڜ>�c��{yX��9"�w�H��g�o�ݡ�J�U�3��v�6$:1��ne
j�.@�H�?M4��;bܸh����0<������y��r&3]z��	ic�Y��H�ͽ�LF�S_�&;�S(�H�쨒��s��+6�oY
M�j�#d���a��(��ȟecs]��2�E}��2/���0|�P.��%�P��Yɭ������i���|�����G�� �l2�7�
�ऊ�|�˭�\Po�QxE�o�b�f�����F�A�7E�&r;�\m~���WQ}1�5*^y��A@fn��͂�Zk��*��fK�i+��u�V�)��w�ln��KG8[��ڛ�G�_-�v�N0<��������7�;���rDߖ�H؃�˛ul�;i��J�vFa2���W���T m�M�Q���%��Y,k�8�ZXF0�r?ɇW�O�6_���"�LR���Oy3�l����G hG�8��g�������yh��V��`���v��O8� ��)v/��I��m�	=�ej�l!�����ҡ����x��\�>�ߴ��7�L���j��*�ȩ͑��5�}Bj�=�ywd{U��Y%=��(	u�C66�����L�������3�2�����w�F�OeD�sW��*D����Ԛ�qg�ғsy��2���8���T�.Vxc�STBi,5����&����i6�?]����t)��ڠ�~FD���ܺ~!���2���8�M����!a�g?�C �f�C��&�����o!����A��j�0'����88u���Je�H�D.���{��j����w"��ɚm�&61�5����м�yF����[��v������8S��;4��O���B��)t����� p8��µ��P�i���v1�����䆑f.j(06���{�w�Y��������Oub>lC�C�	����k��5gN��<��{f����֫�ZFcϾ�C��ii�5`V���F��������,qL ����⹨Ubr1�_��;&
 �J���^l{<���C߁Rд��(7��u�*�r7�mu����L���4W�[4@� �g5�~� _(ӻ4�b ���rL�ϐ����[$������r� �k���9���B)�<��H������w%����������צ���h�f��>2R�l�����g0m�*���| �o�JÝ؅ �˻�]�8s ,��2mH4~�wH�OOA�s(���+���dw9z�
Rj[�F�z�"o��Z��V���;��'�ؘ��I4����؉7}���&���0����m��y�O0�RWD�AeW3|��Q��s&X^��T�1hJ�ɾ
�D��AOyπ��L�h�l���TZ����_�0Qu���[����T4�I�����M�I��B`ymm�b�g ����۶�=���[�m@��	�
=���~��?�1��p��9GRȹ,����Z�b.��1����3�5��9�Y��`�M�ܡ����ҫ�l�כ�AՊ��ؤV$Y��x����y�22����F�����ޥ$�{��8�Ǐ"���M�}R*����wU��^���.��f\w�"�D���K���:�
3g���cM[7V {6�'W��Ў��߫Y�3`��2MYrV9�dMs��w9���ޖ��V�5�O
���f����ޱ©�Io�Q)y�eW.�涅9��2S>��K�
.5;��������K�ݡJ��1ԣ��L�z_����>6�#�$�~���T���a���<ri� ov����:^1�wX""-�E����e3TՃ�V��FH�<�5e`]plYʲ�U_a|��_���˴�[�s�ۼl�:�TXSߴ$�O8��H�k�rc<��E��]�
K�B�1�@UH���m�[Xec1�d%�跋����MGg��g�/v��E	��D�z/��W,4"�D%zK�=��!��]���ReU\�HO�1�X"mBP��M���t˒����#Gec�G���"sX���o$���-7jKnk�o1�ss�����7�V��H��a�}X.�+R�wxR?���[�^�!��F�p��oޖ�L��J�z:y�:���̈�1�N܍Z�/~ �2�.M��[���/�By_E��xv���8��L�+}4�Ғ��:X}��^k�Gx'���[~PW��������eh|3�F�f���8 ;�>*kE��i���'�����1�㐬u��&/�.s�����YX7��]��KF������g,08���G���3�X�*��9.�+$D^R)J���x������TB�ɪ��-m�-
�VF2������<�-�Մ����>)�Q�'�`�;J���T��p>F['YOH�}�E��eO���Γ����À��*`^7C�A+f|�����Ut���*Ze�˓ۥ�:���e{��!zČ>�,M�NP��m}�@����0��{�6^�)(^ud��MP^�*߭�DΔ�z��y��*�a�j�~�H~��@E�_�ӆۑ�| {m�즘	�~���X�F�	;(K���:���ԩ.`X��ÝA�m�Dt�3j�2�M��3!hd���}ynsPςj���4%�{��Vv��}�/�=*��)��ű�a����F�}�?�?ȔK���\M��A�B3���$[�J�̦��&{��y\��̰�!P��M�8�
�2�ϐ��[��.]6�����@�F��{��{=1����/jߴ%lQ##8�.:��x�{I�(o�$��%$p�x��l��Q�r�Ա���J~b��7����- )��r/׮�x����MG������5d�f�eI�e~�JG�̭�C��M��cL�Z��b-��._��n��(�t���H�	���O�����0&�@�;���zH�}'�Q8����2!�׳�6t��WY�45�r�+��7ǲF:Q�^�4�)�5�Qy����(��i"O|�Q�k��jr<���3�����;&?M�'�|��X��ݥL���_�1h�P�i2�Usg�� �mɉE�2ޥ�`X˳�,ڙ��U�;�n�D��^ g˘w���S�M�'��@x��B��Z�|�`
�I��ſ&��{-��ۺE�<�9,E��ݹ��* �5 r�Jy�\ĉ�7Oiy�\�q��_��䰯Y��%��h$|��G}C��K����@��4)TVͣ�K��^m<��oP]�5��X�'C�0_ޞ�Ӯ*	�h0�J�,S�^D0��������R��C(��-U���W8UT�hL�{=t�}h}�~wo�	���� �����W�W]�R�㦈�	W���3RW��_:A+�$i�M�;C�"Z��$R�zUï?���OC�����!��B͢��9TDn+�F�(�4ʿ�qw�PĿZug+?�N���T��.}F�Tְ삋�+�먕;����u���4/Ǻa�|$���yD>}�s�bG�y�1%uE���kZ��1z��_��'n&�/��a��� ^)��5j�l"�hi_�-��v��	u_5�K���YN��;g��>"v�/��V��8�`���&�
}ӛS�g*:%R�@.0-8����F��<�V:H�;�\tS���0V�*زA>l��s�R{ �eţH�xgsȰ�	��ڇ�
,�Gd�<��4ye"�{|��۞|����)/J��c�}s<��,��Zl2�Z�X�D���g��a����,��(@�,�~�`W瞌�D�K+c/@PT���t/M>�t��z%�.@ΐ	.n���yOh�Uk���Y�VV�9[g|����PJ"	����_f"מ��7,�8{��:8|_=�W�A���JRƧ�s�٧����c{9�!��> @ �\�)�C����d�]���?χșصO�#��~W�À��\���H<�AJ���-:q�'�ŏWyTz�O�VCgY
h�q4�A�R{��5?�]��ރ�]Є��T`�j����pNV�2ql;�J�P�:!;���Wi���u~�ƹ��~���y�_"<r��{��h����#�&ۅ�!��e���4���i(�Z*M�b�|�&> [�'P]xɼ�%��z�Nv�{�����֙��`a�z'����y�uz�2��37zf�7V�	�	��<)N;��]A��U�r�u���v[�����h&-���@����r��ӟ��x0|o�gg���?ഊ0_f����8��߆�u���|I�!�V�K�^��)��dye�zqM:����D�֋L�t����9������7�"Ɏ���24Q_�r��%c�x����sTq��U}l��=4r< 7��`��M�ct(��Z�:�p��pQ8ŵ��ܗ��O��zJI����-(Z���B���5� �PTwe����R��A���]d���������</��Ʊ�vUO��Z��A��'.s��)�+�����	��Z"�Hb��z�7�/􃑩��>;C�]�lio�f G����r�P���-���Î�"��]�ҿ��>���������7�0S�O�ǭ\�%"٪�?���C˦뀜��@�l4Cb~вB���E��D�&tקg�b�X�<�-�Ǚ0�F�-@���c�.�C�v�r��a�
�{�ت��Wt]N��ٲC,�)��b?�/,��o�,d2������.�nA���n�n]���.������_��rU /&*��\�����w�NI���c�Zk���	��kw����7Yd�jiO#�Y؊�+t���A�[6��0r�	�?�n�g�������z"����/�����t�M�u%OX)�e ���_�hU�����W�����huGM��R/O2� �hN�	�]��z 1�L&'����ǆ�4�?� ƶ��_�얶��� w:y
]�ɦ}��G��c�=�xTP|�������cDܶ0�@�WI��K[E�g9�d}�gΓ!��&�'�u�4����+`*z�3;3.��V���}d��z�f	�����
��ne�A������a2�ٖ���0%V��Fa*�	�� N�#��`w+ r˪d�_W�Jc��;�:3q>���_Z�IN�I��I�38�Rb�-�ݑ^���0��)J�[�=��J�4�L�1����,�2�oxg]&��c�4��#i�|��2�-0��p}�[o�����w�.�V����
�.Q뵐Y-L+��2���o�m��)@?tF_��Pɛ��' ��ډ�-�{���+X)�I��62z�ʪ"�����)�t .(h���o�u#�&Ú,�ƥ�o����8�Ee$2`q�`n���*h�z����5M��}.,���sڑ�5v]r��t�4������Ә��3�Lcu�>�XJ�mc���7×��_��)}>PS]T
���_�AyY,�o����Iܘ �S25M"J�a�P�i0�8 '7�@���nʻ!��f)G`%6���{!���?yDc����֨)��x�)����	G���!ʅ#l΄*�R��}���Y���y������X݆�4c?�cY�(;۔�¦Y�H��C�S���(颥�,]�?�J\	�v��o��F�;���
���$��EL
3���C#c��9~T��k՞��Kwv��:p��Q��� s��N>�F�OΣdZB�+}�j�-�%�:�T�̺�۷HTV��l���A�mTR�vZ��.��R�<�4{��*8	"�L?||���Q�^�UZ+��1�cp�+�NG���K�N��b,��%�G���T���8�4��d|���
�0�y(�$�r뫅��E$�*"��֪m�b��2�G �צ	��E�y���#�	�A!��c,���,I�O�;x��߈�@EK��r7��2�5A�6C^���Z`���Ҋ�7/y@�
�08�~�֎j��"}tֈ��,K<��&՛�L#$����ÿ��G�!e���N'X�Վ?�Iux���e���N�nP�HE3N�r��w��Яo;��X���o�w�,�I��#<`�6؟/���1]�fW��t��n�o�5v��Nb>��UT�Hb�IE�/�[4@A3>���Ӣ��aה|��E/T1��mI�XM�h�$:��}-TɈ� 2�B���|��Q�wBSC ���.�0�����h�aU�2pLE8����jo5ږO��ID�k�]�͕���8mD���O�
8���gL�2�\wn�<����=���p���p�%-��b�B�g�\,���y�����Am�e��
CBٳό�˙ܶ6��\x�n��qi��������zS��q��͖�Ȍ�;�H�a�8:�i���P�4Y�#pP�+
�/$C����i�W>_Yl�s`02���N��i#���G�NaZ����+��C�<z�=��|y���E5X�_]����&��#Ḋ*��pG�����R�W\�8�����?�R�\M|�%�!�TS7���8r*)��+�ƽ{�0�ȼťCTTi�Tn��J�֭�l��¹ݪ���6ߕ�����N�y�Y�ئP�W�_�$Ɵ�f�xD��Xِ�R�W�	3��H�q�_/��\��S+��	�.l:�
T����!@�2�L+�GYˢ�A��+�ga?��Ѽ�q����fk8�+���D��l�q���*�E|�lT�e����	���&��Li�D �&�M�kz�&pq��Ƕ�q��ь�Ӵl��� HH{Ul��3����IǝΈM�(�V����ϙ%�I�ΝW�����,ES� �+2[��a�F���lI��,'q�/)'��tn�3���p<Wq���e �w�Q*p?��0����&_��*�)e��@H2�*���[mh'���́��?�|�� �"� N41<#�^<S�7���&�dA���Ff&7~�$�XCZ'��t/>�Z���y�=r"�i�<K� ��;^H��$�;p��u!=
d���ֵ����-�qH�ܛj���e�=�ʶĬ>Ÿ�H��j=�M��#�;q)[�LJ���vdPe��%>�nk�r� �3?�����I���.�����{-�!ޯ*=D��43y��Ë���`/��u�Kg�x����9������c�(�I]�A��o8�s��X^$�Lu��+��PL�"
WL͆G1�2'��Q(T�~�j��5�九�l�`8�D>#���h��^�!'Z�	�0���O+D�-;ۦxHR�Z��䡲� �׫����?���[�;��,���_�x
����|�L}$�E�K<�o��,F���&Ç�I����~͜��\�Ѷi�ׂt"w�0F[b�^q��<`q[t�{h@e��/�7��v/zA����x��UY&Qg&��j4/���!��Y:�=Z���0JZ��q���
�?/�L�����U%5a�	�ODnÎCD�CŽo]xM�|����X�5��p�A���4PR~k�a�m�n��jzP��Tٺ+�<PA(B�������l�+�rw�� _
DXnn?<w��Ȕ�ǆ� 8��)���$\)��9
��I�C���	��@1ɴj$m;����`L��2�au/�흉��J�Stc�~�����:k���E�^pi.��=��?�L#�h�NW!~p�i)�G+08f8ПS�9�_.��L�������O����L�z�UȤP"gNEe�N�ԥ�'G�-��Ʌ��@&udsyP�D+�[F�zP��ǂ+g���oš���!�����H�Qx�&P����pv�r�hkxؠmݻ�D�(�V�5K�7^h"*Pʜb!�zI�&�Q����(ޕќ� �V�c�Z���zf1�)��t�1����	��8���*u?'�e�r��4y��/���������K��y!����t��c�r��Ѱ�N�o#]P�Q2�z�Q�;�.�:�8iD�O"��Ѐ)O~�2�k��a���5���'�=��������G�ڑT����=�IݐA���g����h)8�z�6AOv��k*<��j�&>�E.[t�8R����!���(z�1���U����wS�x�pZ%�2�丑�����>��*�[���(�_����#FY��|Q�*S[��,Ex%wg60a>�*ύyR�BH��N�YW{��Ϩ���P-�=���{�����ŉaT�L+�v`h����B0f6�0�z7��3CY��7.)���]����2�_���_����G㵣6Яl�Vw�'��<�w��K�`Zg��<����h ��,L�}a��N:���l���������^ﴆy8Oo��� � �a��^�Fwf�(�y���;34Į,0.�1^����_��ˏ�ޤ��)M�_p�W}J�c)Sg��t� �xٯm/�����Vh1�3_���X;�|�9/�A��A��<k����E��A`\�84&ih�q$)�=Ak��7�I��#y_������M煢a9oe�6���Z�o(�'�_�P]U�R6�W��u�� PC0IA1]N��Oت8E��k�*��op�!}�_T&V6@*���NԗMi��$����,�q1�ѓ�h�PA������`�/���\I	��
����E^����zq�Ȟ'�ۿ�l��^���ugKS E[�{������/�~h��g�7� q�]�h�p��Dd��]������u��*�M��x#�%�}=֌:�$b�E,G�&a�2ʥ?�=��D�J)1��e���&�&y��&ْ�7J��� t�G����H(�FJ#���FDxo���ݭH�H|Ͼ��i�\ -D�%�ܜ���z��"-�k�Mٍ�ｻ���%�ڌ����n
@LJ?�Vź���,�m��˹Rd��;��	c��.�HHnN/��k����1�Vn�XNLV��bM9�N y�I���	��	]m�	���p�#�
u�W�������8r��!{��"�k�ͅ�<r��7���W:?e^��/���M��%ft8�¦����N�Y-�#���Ш7Y��А�����g��i#���~nrbwL�i��b���>�� i�2�"R,q֋"�z�ͬ塴֊oQa��C�4}��M|�6�/��up���E�7"�qw��-�E���·neG��03f&��(eEq�-fL���)).����v<�2a� pH��ɎJY�U��u�^]i���̺Uh^I뾽!�L�'3g�~ROpR��>��d N@�νA�{񫖤ӟ�U�g=g� +�m��8����ȩ�f4�3�M����[��c�|�OI![����[-��m�?�&�ɬ/�q@Q���L=��
 #<�,
�x<1� n��^4}��Ԥ3�
 ��9)�Y�L|�_y�OrQFO��űQ	�\�+��-a�_�LUi5EW�T�����^s)�B���e&EK+�����ҤH�τc���h&-�Z�=iz�Cm�H�V̉��A�*T���������/�匉�t?C�+��}��8���VS���8�<t��8�(l�=����mCcT�1�,�F��"�Y*O�Ni�䥍���6�YA.� h�l��0_���A��n��.6T�ux#�,�������x�{�"���ѻ��a�R:�GQ�v!�Dt
�$��������O[�+�M�"�o�W}}�Wܵ���-^�V�v�&��r>~���#��78Ɖ&�hIS=��{����D��~g�r`�t�*�pf1�i��$�����(�AV^!��w��<���T�#�"5�c8�Ė7q�o��Y�1̀M�y>xO�A��'Z���U&��mCE��ң�+4^y����tUB˗B�:T��w�b
*W�ңYV���_��[\��������s��O�L_j?!O���x�	TV��F��а 榐݇ˌ��kH�N�p7���F��:���l��[�讜��8�_Ȑ�LZ�w�.�}�<���о��B��6�A?��ĕ�ځ`�dH_G1k?�-��nк�������z܂�|ߑ ��M]���x,��7��bw��9�`K�G���%�G��&A��A7#����9�7�{�t�!F���a6�g�:�u���/�]5Q���K�|ZOl7��Uh�1"��,q����j�$��K���e��3�vƲ�j��ev#Sٰ3L��=�c$ǦS"��ߪ��<�Q�H�n]�T��>l���:�Ra�y���J�r��&���[���k%��p�Ya�k9���> �P��u,�~���:b�{̽��"Z�7�<�d$]���:�	�9$�@e7�1)�����M��,��+�t��Gʏą;�\���V�_�A*F��t]uC���L=�X
���O� �=e0c'/C��E�b��yT<�+(1��r[��0Y,�5�'�;�������Hd����{a]�-P׹1����P�3������䵓D��y=d��`��~�ʜ���W�d��ץ��"��԰-mآ����%Y�T�����?��0W����Y�-�Tb<e1�䪓��cT��<���C�����m���>P#Jœ����|�x��� ����&�g�`���Cqp��h>�%I����cE�$��n��U����C�����e!�<��.�I�C��
����xt�;�6A� ��!�̛|�ȳ֜�繪��ú����5�*�-cFd6o��x��D�B�
l���[L��
e���Zj�X�@��&���h�$�w(~{ɮŐ�.���⣙>{��2+��Ʊz+�:Dy�� d]��x[�Bk��Čb���GNAm�A����=V-;,k&�=���T���f��4�	vl�H9X-��?&�:sm89��e
zM]Q����v$uO[4-Ma[�"����O�,P��N�(X�I|R
�ɪv�I6�U��42�/�˧A�+#�ʃ|%&l�лf���4�	ٖ�1���g�[[}X��
��^0�W�qi֩�@��j� tzZKLY�V\{wf/�˫>q�B���Pw7����W�u�����#FC������C�OWJ�0nR9���� ���n?�HI9�M�������,�\ZAൎ�_qz���Yt�E;zM��vCr�z��Ϥv����;on��;��`�|�<��1{`�_�_+�s�>��ꇆ�|�}���(�ɺ�}���Q{�%3o�Nj�D��bRWa����ufM��F"�=>�Ō
f��`v�dt=�H�4�K��iU��䒮(8����G"O�l�t���pGU�>�������z���sI���Ov���1�co(���@�s��n��L�";,R��I{҆��7b�c�r��*icF��g�N<~ֶ�qD�!�|R�9��u��gy�K��ςy�>1��0�ycc�9�f`�yx�xI<�%�����G��`��q�u�YK��+�Q=k���;xA���#uB/X����w���<�
B!(VY/�#Oz<�c�4�è�������sS�<���F%w�mɨ����c�:�	.����+X4Ʊ�`:��9rC�,����[�X篜�B�m�9e��4����-�|�c_.���Dy�-�8r��It�Wr@E**�B
�%d�zM�L,j��8L���A��Π>�Uhz�{BUz�1�M֒�1����"�f��i?(����%���D��甍^�âR�~�㩣�ټ.
^dq��if�r|X��B(~�{���}�扆O�b������%�V��k|���VtxX�_X>�st�5�|�̹gϢ���	w�|���h[���ѧJG?^�ݷA���_O/��F�Vbz���,��-p��= ����h��>e�{~�,�%n�q���=��)Nؕ\���u~�uB�'{�1>p��g����IG3�����?a�뚍��?k���JJ�7*���q��x��*E!��ֶ������M��o�u��(���ߏs����%�"G&OxI����VÄ[oo�Ԑ�<���F|�g�,9V)*ں�ɨ,�c���(.֞h��/r@�����~���j�j�p򽑜L�J���g���Ɋ�sD�Ub1S����}o����>B�>~w��nzssuMH�l�^���$�܏@쒾NN��&�o걤��X�,C��V�0Y�0�L5��=��ѺdbqW�l*���̝#�K�	�xE���l�2 DK�?�����W�G!_dA.��H��Ob/ڼ�o&W�Z�6�M_Z'L�599�Ci��9���':�<��ɿ%�d���`c� �O0�\ă�����q�#R�m��>H�&梢��]<��o�`����ҥ�C�E_�UmRW�����g��O��>��dF ��i|��E�i���v/��gJ����i��<�M)Z�� ��z�3��fps��Xa�6n��nJȣq��"m-r���fH��6-���c��/�h9������������ݲv��H�F$"��i��;����^�%�S�в#G@0�j�q�dH�{�����($�~��m~�A��vY�[�@F�[��:<h�AՇ��P��l�[�/�\�}�+Ҍh�OQ�G���Il4���ܦ��*����"M/W�+�g2��}�<�Ӣ������o����~3�Pڨ5�Ӕ��Z�lL�#��5��@#���|��B�;;_���F�d�I*�mB�pJ���zv	C�H�M.g��1�C�� ��>,�צo�qɣ�1����l���n�Ӟ1���T.M�`�km��`P�ob��,��t�S��6�f �$C��0M��~�4n	����W�����Y��-W_�Kۨco
� wp�nD�]�����M)V�.d�%'m�h�vP��(����U���h+yN�E�����E���	���[�z`�������~y��'�SѮ�!Z���
��/F�C�����GՉ���уCO�����:3yq2�U�"�!6��̨���3N-Q�6>I�i:�s�{h�|�����,p��.dm�O��ե���ˤ0�]�/S'�����%�82|�8��5N��uD`��h�)����n�k]I��?j������A�]���U4w�(^�<˃^�|���.�FPVF���ꖮ���`��⛶�A�0ԣ��Z}6��u�҇o��o�)������/��c ���;$�"���t��{~:p5�8&17���'*�=�оU��5�j7(��A���G����E��\s�\e#���Q%ږ��obkbɋ~�N�t9�»CA)b��{2��k�&����sx.F����-��뫆�|ͧ��Ws�鐇��S}~�߾��	�&�3�{j�2dIl�p8gji�B�u��7�P�wmK����e2�p�i�U��E�Yr�H~�x�.�ʠ��K���T(��#^p+�#ݦ��~C��O�}$��)0|9驴�!�x1���Q,�g������,z=�+ViqS�_mKb@�Y�܄�&uF��g���ݱ��}ak$����G!O�RIV��yw�����KW�n��&�.+^�̥S%�W�3҇\~KyR��8�@�㊟l�e	�d��x+�sLG�N���o�q�����Q���5����34�Q��ӯ�bLS`�����r�b��7�X���l����X�|"���,gM��
�� ��x)��⼠�2V�&��Շ'�=1���^%���[oP�i�	�.?�RWP��&i	Y\����邊K0�8;��$%�e�_;|��<��0�#�o�E��P�H��mK���xt�2��o�iT��8�z���ꉸ
S�*CM@���!���?��p�J��2sM��[`O����(� �����{1�˟��4wE��f��;�q��q!-�Y�ecW�" �+�2\�VA��ʇp륰��ҩ��14�h��+�iY��#P��ick⏿! �����܂ 4�s�?CF�:&�4���4�6u!��;��To>F��5$A�`�_��s$9��s����!~ =k�����P>"���V�-�R��y�߬��x-pp�Բ��eZ��F~Y]��Xw���MƙdS.!H�&e� ��=�Y y�s�)nR�>u� ��+s@O=;��nI�o�u�����Dq-[V+
q�������,��SbЎr�㰽���2�U7��;Z$�s��9NHS>�A�2i�b�A+��X�Q�����9�����:�'#�+�Q,?�mX��ǤV�7�)��$��p�����A�]����;���M�����R|�̈b|�b�����m΁���)7f� àƁ��З�9�8��ǀ��WΑ���)[BД�~�Dآ�_��/C�W�Lr���O<1沎 ���V=Pl�VH۔���R/|�籎���G�ի$���+���5��������܎��M��X*�D����
C�_8��T�9g`n����ɕ����bA���`���V����P�����zkc���/��9k)"[�PӮ�:~��RٖO���+��~+���GjsW��9gJ�1�%�M����W��"�a�'!�<mؑǮ[�Q���H�?���|/�����$���"�P�.aY���gQa�ϥD�� W�u��f^����2b��K|$�Z��xC��~��:��:��߆]
o��;���%����cۭp��} �a&�( _ ́�1R����B��ɔ��'�q|�p^�-��A1:?50�k�B��}��S-,�o���<[�p
[}�䩂o?��4fJ��B�T�&�/O@���W��V���/$C�5�
��az��e+/�<U�.$m���&����������_�=^Ӷ6��老�)��N�ˆ�+u�@��a[�{;c2�0���X��;��*"���Ě�t���~p�i��@ CB���,�F�`����iԦEHe��k��|rشq��U�*�V1b��C�̎Xy��D�|�j �5Է��;�aC�u9�>sA�2�|-V��íL�錮�C����]�2��3:�@{���<�?ob3��	��ؾm�A�����(� 5!6����	���,n�&EN�8�8���=�!R�_�j}�� ?2�@p�M�BN�Iй7n$:���.�7�m�[2���fG�ui��l��R����c��u�M�:W4w���u`��4�Jb�Vڦ���
<k�k���yUЀdTb��A�MX�v�1_72E	������@p���{ПLG��E���_Yeɹf<�Es^��QM�]
A;a�]�y��A�D�)R��#�z$����/�S��Gd�� ��J�e�h䪪b��LH�l[Vg���1�V-�=O�坴z@仲�Z"�?E[u��o<V
Nk4�ڪ��[BT�n:�N��,Ӕݦ�2j1��2o0RS:D�(t<y��{I?��1~��6,��C4���
2^;s�%�z�=R����-/n�w^J3�Ld��0�����4R�
D"Ir���k.e���"��.�	b�Vn)nf	/����<�ê-8`Cxk):ݯl��I���D'�H��t�'x�Xۊ-嵽�����������gW��+���)`c�u�%��[���C��٠"�ȏI�e�U+ArQ����p�i��$(�:�x���B�n�!wa���[P��oR��=L���.I��a��t��]��z]N$�:{:�����E�R�s����1:z��ɆM�݌�*�	��l�Ƌ�hh�3�8��9�A��]�5/��]S��_�zcFW`��^�W�6�.�v�Kf�'��
`Q��f����5Sɵژ~�׆�E�L#�dSQ迶��!�w��N�J~D��U!v9'�ph�%��֟��1�����U������W�3O��:��Z���o`���:��g�0���;4y�<�.�(���_჻=�P�P��Pt��¬�'�q��v���ϥ�7��x-�����Jgش��/���d��Ls,�H��d���9x,����3�|�H<v�Y�Y+l/bVw�FH'q�D�b�u�N)oqL�{qJU���خU��* ��`!ILnd-u�=Ty������q2
D�ty6����IbH˴��h�#��Е:u���g������ߪT�q�P�.�}��n����(�mq�O7ǥb�MIf�7�yX����� ��Ÿ�r���n�[Z�n%�(�4_�}�Y����|��56�!���B����q
Eub	'{�p�mM��^��n��.֛/�K,NG�It��umi�w����tz�C��D�'S��J]ֻS)���7�A��A0\�<5v��P!��r��zm�tA!,HtI�)�Z�B}��T$���|HU�3�4~o��f.��������u�l�jچt&g�P?f�5F�>�\���|t�A<9a"�N�<�a��]|�#T����B��v��#ܝ0��Xdc�A�a�遷�����̵�r/���bd�Kg$�%rD[��B�y<��1�������숍�Jw����Uc#b�0G[ĕ�r�l�����GI�f�����n�����}C��=6Qܱz����_A>��H"��HQ%����ia^��lq�%�k�n-�$E3i�d��[ĮL?� ���ju��25��A)���(%�B��	�}W8��'��R����'ϗt��8���l.8hZ�o��w��A�ΐ$�ȍ�/��@�S��5�Hr0S_w��8�N����~�gP���p�j�axho��*L����Z��yb
$���8����r虾�p�����K��^��m�l-�L�����]pQi�F�`]�(��b���ڡȍ���$�W0{����B��.��G�&��'Vj+Wc�|���K��~�;#IN�V��]�x�Ǎ�\Uble+T��S1�,�U���S®~��i-� ��Q.�5��s?���-'�7���k��$�-����&��	Κغ�'�4�h�����g������o2 i8W��3�C�k^��e��1�;��a3�Ώ�4���,+|$��y�\K�XJ�}wP"��,���/@�
cüd����;[�1j���xy������	�#t���7��ރ���������Ǽ�p��ܰ��L�ս��@��Hb��m�V���(C7 ��6�%詖���
zΔ�N���1E툋��9�%�o�Rw��̒��Ptx��R���p���Bs~<�{٤�I���t��r��W���P0	h/��	=O�ɝ�.��Fq�"$�B�Y	r�ڹG�\�9��_���W�&�w}�a���������a���3��o]�'�W�BY����sb:�O���[|_kPu!�Ii�(E$쏛}R�	�V<�Bb07�����S�t�x���23k.���?�Z<E-�[Ĕ} �҃�g��X$�pbY�=� �_o��I-ao"?��	�3�WG��H �+o?�X��,c�o���If�3/�r����tÉR�"��܈��>���=�E�l�/ee��sQ�ͫ������f�X<"��C�C�'5��iN
�P�qh� �M����O>�R%��SEs �$��a�;���ia�	7؄�ޙ���Q1 �k��v�#�,@{ڡ�/���l���@���sm_<������K�E�c-���cн�����0=�1��KU���������o�E>���t|�|�s+�'�gi���@�3�gq�Z7�1�A%!��HX�7�>_��`W���7>���71�z�5�I��Ɠ��/�<��u�%����DE]Q���-���*�߬�ӳ�~E���#0����
�-"���*�e�<x>7��2
nk�JRW�uV8P� ��R\��&#�
xD<[ֻb\\R-�k2\_0�fa�R��H�ڛo���S2\m5)1�s��z�������;]�����DY1�dI�V��5-������Z`�-�k{�s�O)�xt��z-�Z�C�1�e�Ky���~
}��4�ȇ�%���B�����p�B����\&�����;�u	8ׅG1�/w]����/.��۽�C�܁��LU�l�>l�P#MF��v��ym����˃�;����(����˕i����������t��_�^R
̾��7��N���!�zSpL8�N�l� ��}[4eo�;�u�g��R�׋�|y�Лݴ^v�Y�a�R�t?������r{�ӹ��CR:!R�<|�Z�2� ��}�i{�j�g�<*��x�3��<إ�p7�_`�Y�PO�ŉ�!�%QG�i�e��S} c<���*�Woc�9��,��$# kL	s�K�?�@%j�D<{{�]�&>��ӛ��-Dg~L�lW��Е⒂���1�j9��Tfr��AT) ��n7ބ�|w[Q�-��SHmF9�z!q&l�<���"ݺX���#����U??rI|����+G~��>�*G�?�)k�'N�"���CM�O�P�,��{�xTpi~*�Ƞ��W��?Dd4/SiB Q���K�wǸ�����w�#H:���
N�Y�\�� ����98W
�!�˱��q��ͭ��Hu,��<N<���_��$lԞt|�7T@Z��(���)��h��=kO���e�H΅�w���̭�ی��o�]�(��B��
��,�9�����H�P�gi���E	���� ��
^�9�g}�3![���g����*]rG��@�C�g暔_j��`��V_�C7 *�7�� ß4̲G�a�a���Ł���̝W�7�i����$�Cيy���E��/�7��D
�Y%�ٔ�f�����QY�ٙ�Y<�fS'?0�u�V'�9���.hV��_,�\1��9�#A��Z�ܦ�|��3t/�߄�Х������)���mt ؊p#	ѭ�5,g��U��I���Ͷ�ڒ�C�__U�
�/?�9�p|���AU���+V��GSGoK	s���(n-�/ޙ/�)VI�4�����=��:��Dg8�۴V6�m��A��fi��Z'��� �K:4�e�o��̙ﱯ+
��ì���ʼa�0�0�6�U�6�p�!�f�Φ���_��4���������d���U=BH��X�+����1P�
���ɼ�K�1�k����Ba>u{_⛸֘���
ؚN�/����F.�9�EA!��Xyخ^�����*?Y���[��7�E4��Ϯ4a�Ƃ5y=9�C��L�Q�~M�]���uS��mhƬ53JAG�6CS�$T�T��e���	���}\fgnsSvCd≃4�q�:�E�)�y�3�PkNf\'�����=H�GG�@�?������[��- ��e5�h":=̝�@�x���b�[nX{�vˋ�L����	uQ��+ic�[xu,�uS�)h�E6�eP��KrR��~���uA3VWnU릚��FlKKZs��늵ILi$�w��ɥ5NֺX���/w[���<�!�#>,�wl/EzX_���|�Y���&ف��d��������C�+�-ٞ�|o~�s�����+J��T�*���ɷ&����7W՗{�@w<x�/������h�p <
��$�
u�h��~��@p.FBgꄘ��a�2��s�}����J-�C��ϝ�οz����-��(#�yW�%���S�ݐ��_Ȕ}��l�"������i�fKn�cT���)���&N�+��o�ԚGjJd���� �~�dqOk��h*f����@�5���f�CXEы������ڇ�L;��s*M̬@��l�����j�,��&б�%��+O�����aK�F��ד͝c�o�"<��}�Nй=o�x��K`�!7��f�BGl�Ӌ6'�0���u�4~�/����4���~�R�g�R�P��YL�gX��OJ�ټ^7�@P�~T���X�zrL+��_%�,�� YV�V~�?�`^��AIG<i`����T?&(@��t�(���]xS�Uh��KQ�[؉��N���2�<���v�(�w/��DZo2��,��ށ%������'�Ø��ᔹ6sx�����Q����VaC���L����K���w���\T����H�=_E��{�|f�JѠ �~l�U�f"LCA�l	Djm[�g�ؚ�9���������x+2@��B�D(�i�®79��_v^��ʰ�#BfYԛ��`.����� U�]䴞[������lE#y��cy�ۈ�``�u��FyE��"�p�|�)�O�1���/B=f��7^�D2+�ɦk��D�j�а�(צּ�e���H-��F%A�#�v�w�Fc���{P��u�"�Ϧ���P�'�-�u�bd�9 ���~o �~�Ƥy�R�ԵZm`�;�ε����1aT*�}=\/C����!}:��L?��j[C/ng�^*���=뾋YzׇQ����Т?U=؛�m�	1�?���8JW{���}���9:�T��E�a�SrE �/ SuHĕ��/%bg�,ճ��b�����\��a����������};gl̲�:ыO�z���,o�V����T�0ݢ4�Z��g����b�>�d�W|��B�x'�>��H{����k	LK���>�Xۀ��x[~Y8��zͫ��^=�\& /�ߎ�����B5Gcj9�b�d}]���R�H�fB2���4�\���fe��D��w��"��WOʴ�U���#Q���<�E3�ׅȪ[DW���J�1�#|�<� OrY�=]���u��4����x�����
�\W%�0�ʕX�;�����[5n�<h����xx��[o�ήSg����B�.��879v�A2DK5���NȀ�G�v�����pm��m��X}�7���c���=rPH�-$��Jf�!���C�'�/w� ��&�- ���!�NgM����/NBT���D�V_l��~�!I��d)�8�3�I>S�]\_M����T�#�Fp�:4���P�#@݃u��6T楗�� �ܬ+����<��:݀�k*N)?��T��=p����#m$wd��إ�0����)�5�
��PG��\n<��1Y;h�{�KnO½�� Ί��Fڏ�Mxy�4�+YL���S^U	�Q�Z w������쯞�����d�K�ލb�>&P�eҢ}]�Y[���!��TY4�Q��Qs$^#��+�;f�[��^p���I�p��V�t�݄�P#��;Oh����?�dc>X˂EF��fՎR��\ئ���5�o��IQ��y�4"ڦ@�bf��Fv��fK25��"�_�iBv�u/���O�x1�E�)[Uua}X��I43��(�/5�٤�J�y��Gg�s��r��g��X!+�M"���*���S%�rN�y�0B�`\���]G��:-��c@�3YKb>P�v�-���3�g�'n"0�,��uY�4Fc�����[�U����N�bϮ�wV(�
\�Z?�d�&0�V�˓�{/�t��O<ѕ"���=T�V$����Ov=�ބ�[.eN)�����V+��mDG�2#�'�sPq[�K���Td�!�O��?#��%%�of���5^�޹j�Z�}&���r��h��p�����nk�^[����)���
����>��O���4����u&J���NHl��L�Q�?eR�h�kET"k0�c�MPb�&u