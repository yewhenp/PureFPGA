`include "ALU.v"
module ALU_tb();

    reg clock, cin;
    reg signed [15:0] A, B;
    reg [3:0] sel;
    wire signed [15: 0] C;
    wire cout, CF, SF, OF, ZF;
    initial begin
        $monitor("A=%d, B=%d, sel=%b, cin=%b;   C=%d, CF=%b, SF=%b, OF=%b, ZF=%b, clock=1",
                    A, B, sel, cin, C, CF, SF, OF, ZF);
        clock = 0;
        $display("+===================================== add =====================================+");
        // two numbers are positive
        #5
        sel = 4'b0000;
        cin = 0;
        A = 32;
        B = 41;
        #10
        A = -32;
        B = 40;
        #10
        A = -40;
        B = 32;
        #10
        A = 40;
        B = -40;
        #10
        A = -12;
        B = -12;
        #10
        A = 32760;
        B = 32765;
        #10
        $display("+===================================== addc =====================================+");
        cin = 1;
        sel = 4'b0001;
        A = 32;
        B = 41;
        #10
        A = -32;
        B = 40;
        #10
        A = -40;
        B = 32;
        #10
        A = 40;
        B = -40;
        #10
        A = -12;
        B = -12;
        #10
        A = 32760;
        B = 32765;
        #10
        $display("+===================================== sub =====================================+");
        sel = 4'b0010;
        A = 32;
        B = 41;
        #10
        A = -32;
        B = 40;
        #10
        A = -40;
        B = 32;
        #10
        A = 40;
        B = -40;
        #10
        A = -12;
        B = -12;
        #10
        A = 32760;
        B = 32765;
        #10
        $display("+===================================== mul =====================================+");
        sel = 4'b0100;
        A = 32;
        B = 41;
        #10
        A = -32;
        B = 40;
        #10
        A = -40;
        B = 32;
        #10
        A = 40;
        B = -40;
        #10
        A = -12;
        B = -12;
        #10
        A = 32760;
        B = 32765;
        #10
        $display("+===================================== and =====================================+");
        sel = 4'b0110;
        A = 1;
        B = 1;
        #10
        A = 0;
        B = 1;
        #10
        A = 10;
        B = 9;
        #10
        $display("+===================================== or =====================================+");
        sel = 4'b0111;
        A = 1;
        B = 1;
        #10
        A = 0;
        B = 1;
        #10
        A = 10;
        B = 9;
        #10
        $display("+===================================== lshift =====================================+");
        sel = 4'b1001;
        A = 1;
        B = 3;
        #10
        A = 2;
        B = 4;
        #10
        $display("+===================================== rshift =====================================+");
        sel = 4'b1010;
        A = 8;
        B = 3;
        #10
        A = 32;
        B = 4;
        #10
        $display("+===================================== not =====================================+");
        sel = 4'b1011;
        A = 8;
        #10
        A = 32;
        #10
        A = -20;
        #10
        $display("+===================================== inc =====================================+");
        sel = 4'b1101;
        A = 8;
        #10
        A = 32;
        #10
        A = -20;
        #10
        $display("+===================================== dec =====================================+");
        sel = 4'b1110;
        A = 8;
        #10
        A = 32;
        #10
        A = -20;
        #10

        $finish();

    end

    alu alu0 (
        .A(A),
        .B(B),
        .ALUSel(sel),
        .CarryIn(cin),
        .clk(clock),
        .ALUOut(C),
        .CarryOut(CF),
        .SignOut(SF),
        .OverflowOut(OF),
        .ZeroOut(ZF)
        );

    always begin
        #5 clock = ~clock;
    end

endmodule