��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ���\::���u����N�T��kj��B�hTRZOfܵ���r��ÐT�'�٧���(D�T���S7���;�S�J:$�'U���J�SE���"�<�xI�f,B_O��Vp��ϯ�`f���S�L_>#�m�3Vn�%p�� ��N�~�s����4��kN6(g�I��݉�V�ǆ��~���0{�#�@�D�����|bC��i0��zྒྷ��U��G��� 8��Y��nBR0�[��/�L�4��.���/K"A���{���_-#�'�Ѐ4�,6�t�M��E�~2��6>�)W�gҲ�6�2���s��xS?�EӾ�1�!�AX�=ގ���j�T{y���
����T�Q�ڬ���7a(Ay�����]��&HA�K1�:�b�4�gS/��'���w�'�K|�@_u.ĥ���v�Xef�f,���EE��q�5��_�$�?.;��C�-�]�H�XM׆)�����[����w@ԥ�;��.C`�90���+W�ݳ�}"\kn.-[�՜�����T��`bA�cT�?Ӯ�}���=�$. J{r����҂"5�CL�n�I��dǊ�+�����g��"�i����X3����y^�{ ��-�<�<���|���c��co�~<��#��4�6���x����ⶾ	?�(�iW�X��g:��Z�ɪۃ��,6�A�?6��%Ts# l��_"�rv���DeF���s5+d�[���Z���{�  �nA�'���qP�]z:��̈́<6�G�t���$���>��r��]�`@(*{�z��÷R����^Ķ�G$$�!P��4��ↃMWN�᭧�#�+��^O�⤊���UW߯;���ƨ�tH^v�^ɺH�w,=�����	��*��>Wj��qh��=�_�w�-˗�E��0ZP�g�h6���Z�VD�������|�0�Q��0a�h[eu
�x�x�	�=@ʖ�ev��2=y%����+J�dKNp'�f�2i�l��X?Y3���ß�T���&?{k_�f͹��С�u_��'��)�����m*�->�!+2g-�qnM�/,�$�Ϩ25+Aڏ�x�*��P�x��&]�H?;,� /�6`a��2�g���e�E��I��+��X��R%%�@��:�F�{�}���h�f���
M�	� 1�ӆG
M�~�U�l3]P��� �O0��Uk�Aڹ��;��)�FcМ9�s5�n=�&�j�+v������PD��T
Y�5�Dx��(�`�����Ma~cل[8ڵ� %�~��TV��.���Žg���t�sce&Q�m��k��Ot.�J���ֈ��\s�K�$㘲i�3cZ�?+6�߸C�¿fk^0�q���d���� #���6K1�Qi��]��M�E���H6B;=P��	��II�'1���s�xtF��'��DfäI�f����w��ҋg��3�x���-��ǀ&K�&k�×�a{���%����ކ���F�1F����%
�K�'���mWI,_G(���'˪B�e�4��uYtO�
2vS�z���ψ��YժI`|�e��)�v'Ƒ_���GJi�PgGϼ�B� �_���%�.^��d 3����ؐK��oB��2`�%�E�:A��B��D<7�e�K��K��.�n�\��SZ��p�T]ݙ�0SdbG�v�]UO̾rdC��Gn�v��c��tm�8h�HtӴ���Ô%�W�'^�p��6��i���"�m� ��Ö�� =R��܎��kA��6Pg
e����a\Ri�,5�C�n�0�%�����֙�� !PN���%uo˃��'w0T�ܕϟP6]������;ym��A�fs
��i�������d��9��g/3�/��B��/o	�A��N�toJ�&�ޞ���V$ϕ]�^5�`Q���(!������΂N�if��͞�౺�}�8eA�������ش�H0��p���F3_?e�
�(�#�k��R_�4����6���1��
�]�QlP��x��ZX"�������:X�6飛U߆���i@`Ac��[.V=��_>5x-�<�G� '���YJ8'a��J��n|��f�T�gd.�K!Y^8�Y��]e�N<��<��6g�f�Bd�m��DD��>����TN�V��'rr����Q��wz� �G+M�uO��؎��tD�'W���&�r���Xi��S�H�j���&��oD������Gٮ���ɳ�"w}���}�
�0Y�z�Q#��,?��U���|�p��������D��Y�GFA+�V�ȏ���'�<]���<������v��ï�I:4�L�7���`Nw�y�_:Y*��`r�A������c ��k������.�db�DKM�O>\�9�n�{�)�(�gޕ�K���8)LC�2P��$�ˁ�d�K��$���=km�l�R�F���v\�#Jf]���N��w�-`�}|sIR*�ۥA�1�{�l�Q�UAs��ٯwK��9�������9U��$͋n)P���4�z���m�@t��f��U�,_^�Y�X�|����K���yp2G�
ĵ�bEL��&��GvwU$� ?�mr<��Le'�F[t��X������ʆ��R^d��w�w T�r�m����8:�YsD�;@�!��  r$�>u���K�ِY&U��A����X����n� �k E� �n�S61LO�LŨ�ah����|?w�AY���_؀�vo��Z]�<�y+@Ϛ�_49ء� ��y��J�qr��e�10L�f#���Y��
M7������4��R����}8q�\#�l!F���NY���h`w �'lx�ƍ�;/����|	P[�iֵ�geV���~�r����3tٗN��[�����!'�"�_�h=E�g�o\�'�s@��C�b���r�q�,=�� :T>��	�� �_3������9vH�C� 0{<~���\�
���AkS���-�s�.��gs3�ў2���'���n�&?���I���vxo�Q�e�v��،6��\�.'Ә�:�)��Y�?�{��e��T�o��ʪ=�ݷ.I����od�vj�{&�O52a�Ii��ZY���?)��U����G�D��#�-���5=I��."��6��a�+P�:�����H�߰�q���1��5$����0��M�2���Q�	3YK�pɽ���S�p�w����2K��C���8-'NFR�����եbmA8N�XM6~����6�r�hrw�m>t��h4�%p��������̖�髐eL�����v��}d�d���/r`L���܊D��b]�u�cP���N������hdcLL�D�J���3"�� x����OY�Vp2��č3�W�

�o\R��׼��0�8�Ś| �� a@�\�P5L'h��?�H�%�Q+����7��｝�� �Δc1F�8�_P^�I�]��W	Rlj��q̊?�c�[04�JTw<Y�$e��A	�{��i��(��f�XW��\�~�Ts�x�U�C�d]�N ^��F!�*�y,/
���y�Yg���\#è�s��F��-N9�{:5��W�rC���� �d*������Nv�|9���2-�i�tg����d+v�����k q�11���j�;��(u�d�6��Zdn�ځ�슎�W
Px�<�$�z7T[�rE�<���"�N��B����D���J�+=�i�M�!��Z��ƍ�]�B��-O���#��1^�F�$��Pѐ�Y²_.��ք�J<��z|/,�'����h��pϪ�� A�V�Z v�f;ȣ��"z	@M:c\3�����簾kZ�6:3����If��z��|��M?4��}~O���ϐCSS����o�[��0���z�@7��䍇��St�G��5\s��7}��@P�v@��cr֟��Z�~�d�E�t �W�B���F���N3qr���������pD����Ӝ	�G���x����� 愋���$+�fWJ�[��_��ǋ})j^�;��Yl='$�z�ľ<0|�ʘup�ظE~�g�f�sXZ�d�onh�c�3��`���0���$bg��e6��*ʉ�N˖I+ U���K���6�*�=��z��+��T*��H9MJ�s�U�o��߰���y�P ��x�v��F]�}g9���7(m2v ��_�nF2ble����������_e�tB_0����"�-��<���S�q�V�2	tU@7�As�1�\�뵟uwP�u!��$�}N�R���75ޑ�%{ބ'n1�[A�L�^As���I�����^�vN�K�)�W�F~����Ɇ��P��$����X���g8u�)��.<��	F�YV��|
 �����0�8�A^��qu��*F' �U�M�)�0IR~��)4_ۣ�U�FS��
i�w�q#fh�ZD;C�<e�%~�B*^�g�z ���
~�K����a�K��YSd��m�ڪE*��8����Tj����x_Sd�Z#��;�rʘ��o��̌Y������
�	���9-̪&�N/I�U/��]c�s��Մ��tS�D�Tu8���C��c����̊�!f�,$$fD��2E��x�^ꔷ5�|ϑB3|iv>�=}m����;�&�c�ٵ���"Od�����|�2go\�iS^m������kF�=!C��CLl�ⷔ�MT���|V���J���C}:�&1)��~g2>�� ,�J���f�O|���c2�N��-.0���A&�i�"��'��}��j�9������H�E�(�`G��%�p��cߥjMRw�������1f��d|�6�@&/�H?��W����2��d7C�����j���v�1=	O[/H�GԲ]li2Ϲ�>�D��
j5qo�b0C/�O�b�; ��m�k늲D�H�~ɣd��|�MG|�Z��a�|��s�1q�c�2�[�_-����h����wRg3��?ℽvYa��ߜ��p��C�Z���Iw�RH�X[3�����,_��/8RR�-;�Bo�`6�(W�=��ńk�m̦:���
0M���H�W��L�6���b3�c�Y�TG���=p6J:t����d���l=>_�Λ$����J�*g;ik���{�yT&���/��d>#T"��_�&�_m㠔�~�%���^m�M�8�M2�*�	�h�mn�p�/�x�n���ϳLT���O�7��)�C�5(��̮P~���AR,�ZvZ�`���ޱ�����N_�߄t9he67�9�ܰq�H��te2uF'jv�A���rL���}!��2Y:��tс=��F ���0)�����oY�J9I� 4�Oc�����4�<�OS>l�CT�
�M!բ���(��W��4+?�������-�,I��+��'�Ή�!�;jgQ���ǻh�s��_�Y`*s[ӄ��!i�lķr����c5����k��s�O�������T�ke�2V���BD3���
�N����m~'�) ��eܮ�`�@r�ڢ�=�P3Up�}nT��c���e��iJ2)k�.�R�NO��Hb;�7s����U��w����DE�Y ug4�/�o�$��5V�[]���P|��؍2�4�����5'GV��P�b�P{91���y�0K&�1$;�3��{_ĸ/`���'ʸ������4���X��%F�y��*}����[\Ⱦ�v�%~nv���F������_��k��H�<��7���{I@j�ԱrZU��$L>��oL:H)Ae�+�A/���8s�S^�7�ٻ�3GUNB�]<�~<�%��F(����W�̻�N�&w�]����Jv0P�c�?�*��
g[>>_2*��t�Q�f�x�.��2�B	�^%W�,�}c�Og≥�}rb����?�uWm$�6�_�Kus�|n
��ZxK�%&jR���$s��8�
���F���]JOH�?I:�c���'��6���.�{"<ϼb@#-����+��Ŏ����gr�F���ۚ��ς���X>�)��Ā��[��O3
R[���g���.��`?�{H�{�]?�Ɗ���G�1^
��	#7���{E�V�s!7�m'f*a{;��w%�p�U6�3��V�������O2�%��Cd��ٍQ-���b��h�&�@K�-j];��
�n}Y.)#���j=����c�����A���\۫S����7�!�}�:Ą�I��g�ɽ@��5w<��p��}�L�����Ȫ���m�5�/J5<��f�{���q���1�e��J��E@�p����m V뇯���bY��j�̴��C�?�.��O"��K�,�M�F,G���Ԗ�l�\�Cs��c�{ Q�s�z'����C���̈́$+C�t/��fs���"���i>�|�J#,R��np\ܳr�;sY2SB��d=x`�����2�{�fzK�zT��՗���M o2��a�oI�o��ڌ�jy:�hy%,$�f�,��ڹ̨�JNC�ٺD��X�w�a�e�����>L�ꅿɱ }{q2�rS�$�"ա�ꁀ)r���v��'�|w�� ��ε�3H���-���D���$�=�E�\����Ӟ�ѧ.�
69�?�=��J�����.?>פV�1���݃Ӓ0Qk�J"�a$7���m��+�;�>����b����q���Y�vd�>H#Yt��, sZ����������Vő�7�Ib�;^�]!�ؗ����.��K��n���)��巫Y����V�� ��؎��<UTMm����P���o�G|��rVR\��7���Z�3�ce���:T�I����/e����I�6pTc�&��85�&rp�9�-����C� ,?s��D@azE~�|C�`LFrI�O�^�Nv5�p����g`F�1�� �6�,j�)~�g��f8Y�na���:�6�_�U���&�J���D���WG��j�{9lTcg������x�c�ǸV����p\m�F�G]�����q������M/gq���8S�g<���h4�5��jW��tw+����>͋�T(�ʃ ��=� �X6��&q̐��4�p����23�g�����{)a�o��Lr����Z�f�1�#5�&�5:
��x���pȭ����K-Vz���}&b��`�s��DC�5t�ݰ��Г~t�?g|���L4ު.n�q<�Z��ٕhϮ��"��:c���[TO5�S@�˂
>��A��Oa�5������%5,,����o%%��m�N�9�FkL��7r��������*QU����9�����]1o��0�Q�)g�t>� Յ�zo��E%�TYE W����P�dDg3:���O�E����8��_=�A��2w���} h�A�?	d+Z=�$��P�k��3�)�׾EО�<�e�1�{j]���m����tT[����}S�A�F\n��{���]�1L�dh�����_ �ϹP#�[���N��_�fu����BH����i�^��#+��8r	o,���:��c#"��j� tj�3���]����2Xx���Ł��R/�/ܧ�/���Ӭ��X���Y�vT��'A�eyD>Bh����ε�%7ֳw�d�t��m[yL��/o"B�P�r
«��i���6�΢�#m��"[/p�ܼ'@(���<8�����S(:��(��1��GΠ�9!N�Q�t0����΁��@��)k�%V1��j2ة����ش[3��R�.M'~e��x���F�|Z��i��&�=^�dL��[����\�.�qF�(>i�wz҉�g�@28��0Ҙ��S�@���@�~v��3ܭ��^S�zG)�LWPZ3y�Ƿ�&�"���[��v�,&Q�JF���S�s�Ó3�?bL.#$*���4��Լ��a7�|����.��XV����)���aB��o����i�i,�@��V?����:Tg�a�ԍ?_�����q7��B5N�k��GY%S�������:��H�$;ۋz�v%��E�h�\z3vl�d�{�3��Rؿ8�L��D��{����M�ɞ���X $��^r�A���M\[��JU���l
c1�"�;�ö�\ }5p����O�j=�!��2�� �Nb��X+�j�N��>7�� �!|9�A`LEFzS'����`�+��z�lC���H�e�T �Z��������S��wZ�QN�0D�:���l�,^\�dztp���l/����<Ç�e�S^�ֹ[QO�ܖ�B�V8ylMl����R�L?Y&�NXQ��c�?���EG�fs��~[�:�FsM�� ��h��!\a��3>��/���-�����aT�y��af0��A��~����o�R���q���*Y&���K���Z���+Z�s��]R�n]��̥�/�!�ڥ�w��W��H��P@���qs��"��E��"��2��FR7�B�؃�NJ��X�;m�Qc��hb���x-��-�.�D����5�?�r:��Km��bQޤ�L��7�ɋ�0��Ǒ� {4G�:�ʤ6�����#��0�H�KV~D4�=?�-�+���\������F�^O�� �� %hg�L��*�P�`L-�pw?E���/H�cS�|�zSh�����w�%�w�Q��8�$�\NB#��bCX�.�u�ؓ-v�������^nɝq�d���;�Yw]�P6o�o������d�э�����VB
��
�Z��4#��o�n�)�s��O�7�S^"a�	�����w�K7t.�$y���qV�-?-Y�B�����r����3�^��E��������((������OÕBS����E����X��[�G�.��+I�}=���L~��n��[�犃������c��G�W�91<�\�~�ҍ3�UY���c�]~��K��t�*ur�5�)0v�l�3��7�,eM,8.PfpQ;�h����k�ӽEf����;^�A���	��4�p;)ү���{˭B<���{�D�oe(!�;��v^�-,0gv�$�l ��{d5aw0Qe[�+����U��3$�//O�>
`Z�.�"��Ӻ��%�[�r�r�iX�%ʎ��[>1}�<�V��=B����m�����O�3)%�\�����c!m/�o�5/bAX��Ӛe�� �Ͷ���QNVI���F��f�V�	N�nX����V�ȍFHs; ����?�2��Lv���@�8�A]/Y^���$�(#�[��H�;ؕ<����̐^*�Yq��� yY��ˢ*��ӣ���	� �i�1׎��̑�a���H) �\���Bڜ�5+duQ#�M��o83Q~�,��l+y�G�q.���)�=���٦�\�ƥ�B�v�|��":9�6��+t���/Ű?�U4;�ل�h�O���ypb�Y�x�_~�~W��K�{�\���Iu�
�-�T�l�nX�����r���K�ϰ�kS��W��Q���)�,V��������e�%�K�*���	=���8Am'��{�~v3J|Z�!�s�d�|2/����n�o&�����M��z�k$oiD�}��D�����
_O��O�|c������6�'�H�|1N���Qr`��A�.)<�������g�4�����V}Y_���ţ5�7�9���oE��"��#���+��M��n��ܰ�I��BC��eY�ݽ ����؇��YL���5"��a�uQ�R���	K� �]l�m4'�^v9�r�1(@)5�xW(��[��=���mM�| ��i��jA̸9`u�[�q����؁��l9,)�
5�?��g jq�W<�;;7��6�=���ރ��옵$B}*� 0nsr��h��X\��6�6@qlqBϏw���1��p���j��U!tx��D����S�f����uP�j��܉}mp^�b�����F�͋u�bc���5*�'"7��0�ExK�Ɣ�Y�Z	�x�z�cNh6}]��S�ڍ�^��&��4|�*ᆱ6�� �&����?V��o��6��Ő�ו9ZU+����D5��☚�"OC�zZ���zԭ^����k�or�Ö�\���ù�@Ð�F��܋�����=���BW$4~�tϼ�)��[O��)�ό�B@p��Ml~��C~�TX��AƣD(��ƭ�#>aAɥt���u�����4�#�,/�1�=�~��py5+��G�m�F����[�evZQ�(vr�L[S�d�O���Q�p�<��*X��3�i�h�,��n�td���X�ү���$s�'+1Q��)!z�<������$����L �m(cV|���1C�
�\��	�z�u�s����^�_���~Ik)�j���,�!8D�q�Ho!QY �0��>�05���8 +���t�8dW�N|�b��?�|�!�2A�{I��p��qiﷸ���Sea����Hױ�3C:Nŷ(�@��?s��!{�0�(Vw]�W�����ϐ���:Ĥ1:1���0�����?�v/s�
,ے��j�U�xQ����c�çb�vd��T(�M��2��YD0�(W�o{�b���?�9�֕b�6$��v��^zߝ��G~�߂�����1��ʞ��<�)A��+��Ύ���,Ϯo7�xU���,��~���Ǉ:3=��1ơ�J���H���4{ՓG/�7�Q�)��ļ:���Xf�YcH��0W𣪢��]iLb�&����/"���
�4�ZgI2jmFDV&�>C�e�Q*OD�2�P=;�xu�aKzM���|�3��v8�CP-%��Kz�`��<�&�(R{E��:��:�|��y���ԃ�\���A�*�y�޻�I���Z�#]z3O��`%�0��z��Wo�u�R6�-�蛭z��:��^�����*?+'�~S�
�D��H�Ϲ�9wLYʕtV�m��z�'�;�T�:||��P�:��7���jastC��K�sw�P���	�u�o��S#�(���Y�-m6�XD���V�ؙM��֪�lC��ב��P>��%��W�o6�N�{)�����bd�34�KWWϒk�>�LE2&���S��Ⱥ��S��K��hG��gF�J/:�Ξ�-3�e��;��u)�R21m�D�����6x��9�/��o?��������6����##�����8��l4�n�7b���c޻���;W"zmZJ�H���Bp�����u�~e�SNG=t�!�J	�G>	�����+�*����q��	<�[Q�E�?;7�Zׄ,����Q�#m)��׻�nL�1�آ�`,�>�U�gQ� ��5h��r��+����H7�^W;���ѐ2�V�ㄦ�szH���m��y��R�@�/�n@B��dD�eh+�t
8�u��%�n��D:�o�gx#�Њ9�+9�K�F)�O#�c��b�|/%��)�r�(����Z����|�T6H�#AW6�
[G�M�k[­lI$�/{�D;��(i��}l��M#f�!�??(f�r-w����?�����-�Hr�P��cu#rzbň�>L-N�'�6^�u4�-��+��N�Rl���K5S��$#[�2j�]���VG���b�)u6��S�]q�1������˼����ar��n�5r��Mv}�
rձ��v��>j�i��|w<���&�<نӸ&7��A��[���
H�C~8��  ��3��AX��('������ODm.��6B��7����8j�"�^`�q�
��l����OT��U2��b�c���&��\#�B����S�Y�	{��"���q��r���,<7��[s2GTV��D��ج2"�����\���ں�b0���?�6\�ƞ=�`�r���D�������������W�ͪ3��yz���V�̷A��VtU��2~II�>WVT�^Ke�$�hL���a�X؋�������a��%?4�e�����;kE��7�ϣA�d݈v���v�ۭ|�s@=���N���k�ɦ4JgF��V�+��]l���)��2/@si����A`E���J�yQ�%^t�k�|��>�Ũ�a��A-�����Δu�Me;��`^2Z<��G��wZ��XB^��UNV�����X>����,�W�$$ݡ]�YQ��Q�8��%��WЃ�ʑ��l�&��$$Z��309����4]��4������s��4���	¡�@�I{c�d�0.P]�|���g�|9iS�D�a2�Fmף�Z/�k����3������4M�8�m���
��%�ks����H�-N��Å�4!!�Ѩ��#&WFPx�d,�my <��pQ�+��{D��Hݯ"H<y5�����w���;FI*����i�:�~�$�2j���b��V?Ѧ{��������M�Q�Հ��'�*�Z���S77US�?)�Fw.�X]!��e�T�s�a� �^���׵��M�N�,紖��wHP�K��Ţ5	H���(�U��>O��j�yF>����WY�vW�2�دx�X�X�/&��J7S�n�۠!yFJ����F8B4R|��F�������W��DhngW�+� �Ynl�z��;�'�wv?�0qtO8���px2g�]�He������u��+�W {��E�r��q��"��8I}�!��݂���1�ji{c3d��>lcu�ge�0 x���=N�D(�p**�t�~��ֽ��p���'��`�]6JD��(q�t]:��H�%'�}�����|�3�-�M�ڀ��3&_��a!V�41�Z	�ND�k������5me�C
�q"F�m8�ω�:^��y�(x�kTbXO��:ƚ��ͫ}��Zug:�M��G�a�c�QhW��b�|�]���?I�(�q%T���	)�ԋ�ʰ+�Wn�\���ez-�E$f�3&����+d��C��m ����Q�P��~��|c�v��r�qݣ=j�b�)�8(!�*�<�&����ϧ�1@W� }�Zq�͊ua0�W���WhA���>�k��f^Хq?���ݲ�bm�I�᪕��Ì����	��T~�A�sMH �A�b�z�{�U������cز�ė\ݠ�CW �H|3�K�A�s3�)�:<>:��u�au}a�����
=���b��\�T9E���-��r�����d��e�z�٣�Y�����S�� s3�����h���.��ޤ��e��/��A`����'��<��s�<�q6?噂����.D#<�����X��G�����^"�J1�2��c5����$��q%�4�Fm�\*��ϭK���lgN4��a�����	��e	H@/P���(���΍�ktn��&���o�$0�s�b�(��W�ZB���я���p��/b&����]XK8r��!9��k���0�*9l��e����䢕�q�tRQL�e��}�q�΄�wۃ&{�d���y���E�"
�E�֧֠��͕�����,� �r>��5C0 �}�����7An����p�X�2U�a���+&`��M4uT���;̲��u��"�f2�6җf�>���������m\Q�V[~���������d�^���a��Rʁ�+�(�B��c�b���C�:<>u�W9�u�;�P@�-\]�^��Bu��:a����Ȑ��v����>�bmC܆T�����"t���씜�£/Y��L5[;��az�`;��l��o��W*��G��P:(�v�c��V�D�����"��h*&.��\�/עP��M�ߜ	���8�A�<���)z>��V�~i�&}˞ ��G6
�bXʜ� ���j�
u(��Z/{i:�O�eș�G�n���^dR��{�M�w�kL��5Rg�<��}����PА���ھ��ȳ?z=4KDQW��}ϯ��ve�l�N�q�^_.���ֻ�=0��Bu�a���#����zzڠtǫ`��e*A�Vx�0���33���v�"��	Ԃ1�x�����(f����%[��F�o֦�������r3H�hsQ"�LY��}��=9��_� �ɨ�_�r�4��d�L�2��3����%ݑ� N��a"�ڼf��V�����b�RB]������_��Ϙ��7���B0@��,ב ����\Cv� X.�x=���XII/��jqW�t{R�>V�#'$8����vˏ8?�������X��:};e�o��?/���%�����b�e��CYДx5�Ɏ&9ܙ�5�~a� ��L�>WU;hQ{�����SʓPrsCd�u~��V�=��-��e�� ���`��I��m��Õ��Q�0��dX��Q7 R��j��j�`�Ͻ��h�T�����-^H[���#ZD��l��mE�ǧ��](���A���\��}����:l�c�dG�~?z�E�E,d�WԚ���R��=uK��}�,�$��@��i�Sc~��miM�b5��"�lO�b�s1��ϙi����%���������N���mD^*F�f����[#,��VN��9fA%c�7Ȋ`�We��4h4��-V��2�n����o�F�V)jo�9cS2 p)�p",,K`����w��=�z�
B�K�,w(�e�?�u�{�-��^=�v���Z�.x~z�f�)�B����f�,RC��K_!���#��n�(?#]��L���*�W���1`�xc��a;6RڤYc�0H�vɸ��=�ﻥ���4�6*�%H{���+��,�w�����FHn�߀+W�H����:��ט��BER���ƪ����O.�\��x���<�ķ������D�>>(hY����
V 0Z���2`��Z�Q���,r#ܓ��U��oŴ��\�kh�)����Ǉфϴ��t��&w8��s�j��O� ?9Zt�������@�0qM)e�1���Ď�F��	iT���FF�''��i��o�
���,|�!�n��,�@��Zj֤��#���{s���[D�Kc�,�\o�c�pR�����0� SrfF�`������Wl�c1��P�M�v~'C��dE�[��U���t|�Yx�l%/(߃XI"u�ng_�[G>{�r>�r��"���E��%՚��{{�_��)fv�<V�P�t	$I�d�O Έ�B+�����J�2$������/N�Лҙ��r����)����K�.v,s�^"��d�.��1���
�d��[(͆���ĭ]��"i�.�	Փl���&�>�cu��>��9��>���,�Q2UҴ�Ԏ:���)�n�c4�5N�4�d[�Q�7��S�p�E�Bb�&'�p�=���['�$E�g���'ꇾ��YޅUUEm�I��{eOr.�=���A�A��5,��/nPE[��{7�Z�Q,a5�z�#��+���:��e��s �e������E�}�����Z�N2��'�P"���D�S��W��ޭG�`�ӣm*o��p� �������=_;����d`u]#�{H�p���q!̔�Y�,^ݦ��׽�u�Ś?�ےW�X���]�B�����,�w7��aH�񃐘��W?vʸ�'��Ⱑ�z�+�_�} ӷ�z�� �
�����]��(�\��xfn��E��=�U:���^o ]����F�B*���=_�0��P� #A��{$pp���"�=�.�'�6<@	����ң*���:�-��߀�����u���h=zC�cPm�L�Z�^�zn�@\T�}R��