��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� s拊�[υm���|��ק4N��k�I.�=�]cS�����9���Ɂ؏��=P���o�\��!sV�c��|�bO
�(����w����u�n�q;�+�$8S�N�EsB4r��-��o�-{V�!A>ӗWR	���3Ini��2�M����9�
/�ղ�DNU����(k���zw%,���]Km���z�Ǖ4ヺ���N$�]q��ʠ�� ���<�5HtE�uCq�,a���/FM�2b,�R]Ui��ybF���i�'�ݑ��p[MP�����w����{�t ߽�mN�\^�~���w�B���^.�N?HjM�Q���B�p����p��!�i�B�~B�C$��I���'IFI�T��B��U��F�2�2D<ӕ�@���AȽ#�	��j�`��<;P��8Z3�8���_P�a������,�����seK[ u4U�� ��Z^�#P���k�		7��i�(�vf�MԵ�y��ZM���NI��C��rA�%�b�Kla�ʟ�-L!| �Gϛ񂕿�/�}ٴjGv	B���Y���A+I�M{ �S�@Y9VB;t/� ��!/�J��b6���q�N��q�o2z%|���!����.�a�z]Iw���F��$��S_�i�S��un���@��A�<�ݝ�4o�̏��ƴI8>�[��I�S��.4����X�h�2�Y�r�`I��p݄�4D����'�7��jT��*���0"��\���j�}6�X����">�u�D	��3}���A�xP�M(��H��˧����D.m�	�(*�Mbr:g.��ۊ�9OC�15�V.tٕ�rC��eo��p�鍢g�v�Yk؃R�ɜ�+PC���rc=��,�����?s6=ܠG r3�0B�[�����5�Ҥ����Q��ɻv��o�iN�\��n`��W���1��t �E�K��ד�BW��j"k��?��nY\��q�i|#E�����+�R�p�/+Y$J S�g�`fFӵ�NQ뇛_e�%3�w��sLM�Ѭ���u4fQ�_I�*���0���'���ѳ�������r ��wT�:�E��4�A�ý�rK���� ���O,���=��壵쟴�P����;`���n�7�)��.p��:@пT��	Rʋ�p�J2G)��'e��=�&֗�Y������;�����>_�չnE���Ht���Bu�j_@���Q	b
�s����$lӒA^��czcb�>�M�!�K\!��;�t�#�T�o�Ol��ь(k��1�{l����/;�3\��`�<N���i-s��JHp*!�Е�]rq�V=I�i=V�Vd����4k��������k+�c���zN�C�H|�"�8&՗����K��>��s��]bl��1)~"8��$~OF�.��E��Fu�e�>�k$��'`i�@A�Ҥp���IzoWf��T���ț4K�}`���C���vV֙����jr6��=i��s�8��x/��tM(���/(s�%��σ2)���~�*��P\��X�)5c\�oU|F2�?��-+>�����%���=��۞���a//�͉��冔�CHh�x�6���o&!�9So(��;09��f�@[M~a���l|`>���]�#�(�F���k�b����4�H>2=�/��8ڞ�$��PR��F�)�f�q���IN����'
�y�Z�dd��r��&�L�� LV�<]׺�Wkk0�B�Cvi�[��pN�����^�����=<#�|W�W��X��2��?�y�#�-�,�d�l�)}�_�뭴X�G��M����_��2��V��M���#��z��`hR!V���>lZ�_��� I�1�je.����Y�e��Em�Ro�^=@#W��m��映[��«ժM��Յ�{�OT��{@���/�JA{\Vϲ�RT1�c[߼U0-W�Y�����>Cl��k���wEw��,�?���R���_���<�I��I��R�I_���>�*t����C�1e��'rxZ!�R�xA�A�r����#����v�����W]+ʢ������O�(FL����f��9�ް����jA�P������s�y�{����dq2G�uO��Q�bbH|��ZXtibAk!l�ů�q���%Q?/0��Z&���*�0ԋE�J��F���
R�(���)�db�[y�>�6�LW CW�L����0Z?�9f���J�oEU��կ� &{�r�|���H�v�[4��2��e�Lj*�[V�z֫�HJ&4㯑l;��n���aX��s8��� !J"^F�Y ���� �U�3�m�"��F�$�=~�r'�՛��_p�M����+2[�p�!t�g�%��1g�T�0�G6��e�k�H.*�3��*���� ��a�I$��s�tB����P��E�_�1~$��F�6PL��̋!�O��� ��G:�>��6�?�s�����]��g��h7'��M��bъ�K�	�\�E�q�?�3:%��9��$��{si���ƞ	�},Q��;f�^|r�]��gn#���Z�I*}�mf{�������z���-E�ud��2aN�W�8�ZHkH���TS�E|7�a�k�ce�ì����l.,5A�(aU����j�Z��Tˢ�γ2�����>�)���tӖz:t���b�?��pnlTX,;#�u�p/`�&8�k��)�����^�?����A�HZbo~���8�C��Q\�պ���i�H��
�������hYJP�����JO�Ļ"L}�������+n[+��2��=�r���a����0#�����T0�����qE�-V�D�	�%[~�6�Qr��[��9��!��"q�Ԧ��I,�c�A^���j ����.��vJ̏Z2O$�8���V#댚.,�����s���>B��J����{vȺ:J���?�d��͞�ѯP�ͶC�0׷)/P�)<L/.�����P��B��i�ʍ:� `[���'�y�k\{�	3_��g;����}�͙X�����Lc��~�n���?���m�%7&P�|��R�Sd8d�	d�,�b��G�:G�̖u��V��8ޟ�%��Tv٢��s�S]�U�PN4V���BoR��\VYp�k�r�: �ϼ�����-Nˑ c�'"�/v���B���\�.������������e�4'��7�a���)�:{��k˭��?e�i+�B\�3i�^/[̀!��R��-�p�vw����ï���5�U=u	�'�i="�(l�|��|1���1S䛆A�����0d4��(yjMC�r�%�R��
����E���^�F��)e�u"U6D�7�����̎�	�ҍ�k�$w���%��l��<t��h�o: Y���Pm�ߦz$�e�]��8�����#�#�@v�Ӿrk��h���f�<�'��Y]��M�Փl��c�d�ԯ��$���3j����!&����H�J�x�f{&���$ʇ��k7v;�����·��oDds�n�E��fӤ�����Q�)�c����`��FL�+��r�*sgPW?ǓB�hw���q�����W����;��e��?����3��.�ۿ"�ü�6�Q�˷%�8(
��	�޸�9���z������%�l�3�'npsOE��[Tx�x�sey�V�l��� �&d�{s++S(יi��0ǐ��a���ѱ��Z���]bC[����t��O�t���� ]�KN��I{vT�����d��-FJU$g��P�Z��kbP���2�� �%K�k|2/��n/���#'r�Hٜ����Yr��B���W�p�~Q�5j��I��@���A^,A �8��j@k	��1��Lz�%8�t��K"{^r[?Q��Q���>����`("%�ߗ�zi�"�^mi���]L/j��w�S`L/��7G�]ȃA��=N�� ��d*" U��4��6X���9
_&���ꤹ�]���D�%���Y.+v�ty;O�R�V�j�ky,�>�����<�����g�)�J�G�]0�o�.ݢ�����ӥOI�S�҅�^�8%b�;�q&u��x�&���"<Fg��J�0)Ҍc
p���Y���X����)$>�����	�3�D�W^6�3p, ���f�ݲ����I�� ��Ti4a/���w�:���o�vu
Z�@K:Ok.�o��"?�ήTq1�G+�������}D�#`w�,Y�b���P�j�^�^60�� ���t��	e��$bl�[� J�;��Z�.�v#0)�����+^<@U�	��f�z��%���*��:�N����J��?�H��q���n�_�u��UD���Y��+���WLT�	%����C��I����Fg�x�o�vfr?���n�Y�~�^y&2}!��E��A�ci?+3�ԏ�e�e��zn�MU�s6��Oy�,��0��n���،26�G�+ȉ���pG����*_��W�&��k΍���m*���D�d����(�f��Fp��D�ܜ`T͊Ȋ��;��c��QTi�"�WB~9��Fɸ��X��,�=�/�w�8�8=/ �3mn`��6��xw��(-���ӵ.S'�ȋ� A�* �謿[ԧ[v�1,����A���0	�:Wc��D$3��=�p�a0���5���j�k�}�E�4�/�y���َQ�{��q��IB��BDP����&h��o˥H��z���r���=�����n�<ܒ 0�~��HjЎ�h-��e�?j�V�[��ޙ1V)����(�/��Ç�Jѭ�r���oۚ��h��c@l�?������It��O3��#;(4�P!8o�b����a6��4�e��Wѓ_Mo�L[���{��e�)q������`���R�Ii_���7*m����Ʌ�^p�KZ��t�+�ꝛ�o6>���A���$}����Id9��q�J�d��jܴ�6Hs�_��A�`�UG%�R�)�4�&��-�J{ T�Ϋ��ڎr�r�2�*����j�����+�e9'r����S���hk=�W�S�ǬRP۹�2���$�/[u}Ō< ht�s,D�h�Gs��=4�C�h��W���"����{��B ��[̵��b0�%C���5)J� �7��*F_���M�1Z�К!Y��BK��em�'+f�Ƈ�	#^݋���jh9��L��)��[��z��"C�I�ȗ�E��x�S%�Ϯo�S��i&A�������˹��n(8�I�*����p`��$��tb��'xr�.;H2�i� !��qA9^��r�%#�G��E��3��#ī:��d?��o�mk��UU��Ϻs"�EM7�jyD���+����o���>=?����Y�DM�K%�=� D>�Kj	�Q]B ��M���{6Kk���|9�����h���k?�F�>�ѳ����3���w��%��،�ԙ���ȧ+�Z]�H~�Uq�pUvn���*c�q�c�����K!%$�TV��Dv��p������8����W�q(�vS?��-�;��W��T�h�ԑ�~�:}�Q�P������Q��817\70=}6���%�����I�v��vx��fȢ��[�:N�y^BV��D����C��nޤ��� ��B�<��:��ʾ�WRr��A��s�>�����?���8�Z'(��I�!�B:W���Yi���Q� S@C<D�0�f�Q2�R΅Q��NO�W7j�#��T�@�26ES���G2@#*�>��x�?/�U;���yc;�.È���Ȝ�oM��42�@Y�>����!YԞ�	h�a�Q=����^�����W��/�t���{b�x:,��PR�
����[P��oZxAE�ÜS�V�j�r��4�C�'i
�\Dv���1��(�L�f���7��ڰXZ��U�ȋ�<}� �>	f���:��P�
����@���s��s�ּg8��2���FyQh5�\�[��*ق#�����-4.�:�����,ȯs^8��p8��;��Y]m�:*/�v7U�2�����ui�J"6�ֺ�u���L��q4��ވ'�==�&H/� ��k�c��}�`���
��t���{' �O�X���,=7��O�ߘgc��rYc�tV�g�8Zw&�<��pD��ܔ$f�A��|�����n��,�������Иd�4��;c��X�O��mO9���2CWAQ�/��E���ן�	��2�������*~[��"�φ\�O�wH�B���lH6�֎a���k�"��+����l���Q�~\~�X����=6���MJA�z��A Ԇ��zo�#��i�Ί��4��E���_��}�<&��A��Ĉ���1�E)B�3�a�*&�6�~W���Vi��혠���?�	�Z�(q��C��V�Z���
U�$�>|��ښ������J���"m��Mqʴ�Q��eVT�"���ѯ�[4�)�����u��c���4��T~�����h�"��Pr��>"*ON�:(��|�s_�`(�K�Vú��Q����H�ɐ��韮�ͅK�H��N�e;�ۜ+%#~?�4�1S�ې���[^�J��l!�[x7F�� �<��{WUy8�F���~�/�-T@i,,-����YMF�8���^
&p�:Z�xw�V�iT�����PϦ((BfB �=��Î�T�*��얦Վ�,��"�3�m\%��b��@��k�]�E(�\�pnTM놫��g�Q���[�<>�����$V���H۫��S�����\�Ѕrq>�T�
���ph�r`O
���u�ҎKP��n��mN��.�Qd�<�W�ArðK�����"����j�O�%��>�/��$�I^�p?Ϧ4�n�K�ǂǗƷF/���@`[����)� =�u��=5�o$��L`�ţn���~f�VoO�Z`�&|n������l�D��t�kO���4%�3�Ƚk���Hé6��*��~��ܱ1�c7�M��D{�U���@1S@�q��t��f��*�4��fz=>�