��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� R����q�m)9)�L���dh���~�z��>d �럥h�z��Yr��Ѝ�6s�����^e���j]lGI�(V��K���'a�Q39�aUgv�=���憛�������d�<{@��������(��wukt�,���JO���ԓ*�1��ݨW���Ħ"�"�M����|=�� �	"1����y���t8��m�2�
�JR�z!���Q *h�r'*�l��̓�s��0c�ز�ˡF?=z0���ؿ�}@F�fr<] ϊ����_����?c� zv��&���xЛR�7�ɷd9����QToƳ)~|<*"a�D�=<1����W�໫��!�u�; �8�6����f��g}�Rb��R��#%ބ^�L٘$J)S8��H�1��(���ª�|i���	pQ��n���$�R�E�^&�I���a��L���f!�*O�Nwj����!.��g���8��-N�6�qY	�VQ�J6 �p�bu���t�-���&h�i��a�bhIv6����Y�)�~�Nn�<�!��;�I��)3�w�"�����"��e#�2��.�@�4j��3��eX>WnQ��?���1����i9 '8�N��UR^)$x-�{��,�5y��F/4e�~�ܙE��¬.\�L+�]8��+��9'��y�[,�zBaq�BF�W`4�`��
N�顋�L=q����3_�������.W���S����L3>r��^@�B��EV��L-R��߯H����SQ3]&��g�lA�,O�o���}�����EP?�	���ۼ�4L"��N���q}o�!��H5�N�?L�暶*"����e��0],�s��u�,�.Y���{�%�)�?^�sJ �tD_�b���v��/ճӱ��T�,%������S�����9NG7�A�P-�@!���� �Q�j��\�ty�T~l��0I.hgO�����p1cA=G#5�qio?���N�pp`��"�D!'#����Îu�IMړD$g��k���������Zj���so�o������Q�d��j�ў����t�''.I�{0�R����0:��-�D�
l)	2S����@�x[#L�Z���\t��H�p��yDx�Ws��d��z�r�UhUk��&�P5�(hU�Q~j���/�:��e`,MBt�KP��:XaG�ک�	��Mj>c	koDm������ZweZ�
���%ja�
t�zb����H��(�.OtR_�x���p_`�6XI5��"@�/|Fk{i.��n9��宄����xH�_̲�H^�]����bqK�6���d��k�*�?���L��T��5���B����P���i�POw\�S����5���b������X�?���S���#�oH����� ��z%�W��<Eߖ�v�ŧ����~!_�MP��apt;��e.���=1�JuP@|��r��C���hCG�z��	>��,���$E�$C�뛴�g�rxh�G��RA_���&n.�.p���{���Ɵ��T%�	��q���D�U�t�B��R"N�ۙկ�	ޜ��$HeO:��b�<�[9a��}I���_�� �������,<���L=��\�3�A�ֲ�T��u!�O7|���m��K��*�U[ �ʂEK<�P�~j0ۦ����}�܏��q�-4��C�{�m|��]I�X�>y3�@���*��G���dc�{ѝňɑy4[�:�O)����=�x�k��+�N��4�AD-������{?�~��+�<S���ީ�9��9�$T��ȕ��r��)����EF���fio��}�都�^G�Q_�w�h=�	<�T@~����o��h��Z!�t.#���D-,�u�gG@zA|�S��s���F�D�H���jX�ݚ��J��"�z�[��k��zm6�7s˻_�U�<��D��-��ef���5����Q�;����/�nZ۪���aR�#�,'��e��r{���]8W�萶:���Rk`�ӂ����� �mK����b������߿��sl��)��)���V.�ʔ�rTEHߝ|r�$��s_a~�겻��}���]D�J�����:�������⿰�B;��G���p�m<
.
�^�5��f���K2+k������'?*�%'��f��$H��b̫kfa�5c,60r$��*�l	�<\���*Ub�]?�?���#	���e� ��x��"�L���"�Wؽ��_�	�64<��+�׻�&���Tl�x����X
k/�������R؇�1�&�/��-xd'�`?\ h�b�'�|�>�s�	[3��.��精1F]}��(��k��T��3]J�������h���d�I�N��,����T�;[� � x�:(&U)zf���{ٗa�y�d��y<���N���/G�Rx�F��0`��˲
+��&�U�``��{K{!aAs�[��'���h:�@�W(���/��E7U&~ n����0Y(�[��x�������)A��V@��h��C� X"�
u'Zgx�G�%��r�֢��Q��.���L��/�IIs���W��%��N����WF���k)�g�3��x&����"���N;�c���i�'�"q�5cQ��E|㶶��@<�E`�p��5�?�5#��O3�aը�ɱ(%�c˱
����T8����6og^i 2)s" (x�RHa�cO���3�F�Nz��Kc`d��I�����n�ߕc`1hL3�kd~_��k�>0��[)��,�|�=�(;T�$lȼ��ǚ�ŵkͷV��w}m�>Q�0RX����f��J�F��([� @�p�U�#*uo�#o氒#~]��
�J*e=���+�?��$}}{ŕ����3�h��X��r��;����R��ܚ��I�~��i��.8Q��D�s~�L��Wa5��{e1��Q��70�x��((�QhY��TK�X��;�G���)l�|U��,�z?��w��9pUR�x��& K~B�Zae�˘^��0)��:/�]��%�ʅ���n^����<7�Y��g�nr?@=V����P��3��6al�'��Q^�m0A��W�S� i��;H%�\���CR�f�m`Fn73��+���7���.�˩[Ԟ&�'�^�^�;c������螮G|�)"J	��+��� `l;¯p��v��8!O�.,/]��Tef5��ś�L�Y��V3���(�����Ւ�_�N%�I�<�tJ�޺qt�L��B��}�u$v�Y��LY>D���)3S����8M�$���RCO�9�'2�{��S��#�[�PHK�I�o>/񝷖���K��B8�G���>Q5�z𿡎��A��ξ��M�Q��m�����eH}�hD�wDuj���2��B�P�	w��'��"}f�l,��@حJ�g�t�g*�&��d�k��-��w胱l�D^j=@���c��Ń��R� y&�&qP�Ό��/C1���J�؂V�ju�W����M�f������-�W�k���1�������G ���:�ǃ��~�gn��hǕ��s�];h�i��Y0���t�m|ȉu����
iΐg^9Lx�M㳝{k�@6� {��
sl���'���C����	�����ᒄ2�ޣC�����'KnfdG4��Q|)��*[.�^�ͭ��L�A7*ـ1D�������3�������g�3Z��@::b��*q�t^���G�ƕ3���6u��l	f�FhD9� RY�a�5�����6&C�mC�
H/Q�&ܢ{�����j�\BK��N嗾�!{K���b|l���x�Gvlk�k��Ns&K��
��tsE�?���?z0��ƍ�W��;�/�4L�5ڳ1�h�����ݠ�8����!��$����pmPH�N�����+lQ��c�o��/�4ŁE���H��5�@Y%(=�e�� ����$^^�� �Z��������+����D�/�#>�v��.���Q���"��r�]ȣN֍�S�i�#[��[H�CR��yB��؍@B����7�n�%�J.��{3�Ţ&��L{��ؿ3��YA ܼ���V�}�O�ݢؑ�ݦ�[=��%3q�ށ���(ǿ�'���U�N�?��؟�3F�B~���E4�jn%���;45�Ǘ�7�ep��9�Ƿ��x����
��.��Y`��4~N�aqq�����ssq����0�-�Z��%]��M���ue�i�g�j5ku�W�q@t�L�U=G��>������N��� ���E�N��ӧ2�}����F���P��d���"��i�߄��0|W��i'y�ns��-�s��]��e�,�z�V®���U(��a[gj8�hd?���Y���qI�d*��% i֪���lv#�2��\���T��NQu���Ct�|�u��A�z��tr�������2�F��K���B�W�äWӢHȋ��Du�>����$?�9sJ#9{���3��Rs�r��[�ϱ���L�Ou�z�t����~�NH���������]ZP�Y���P��5k�����Νo�W�hXA\���@h��s�T �qJ��{�J�v��=u��_R�y�͒�WC� ���k��GTU��>�K�p]>�d6zm��^X���g��R�Ֆ	�\ێD��q�"�}�kh��x�/�4��7���J'B<ط'	q�p��k�_l�[���l��#�(.H�9A]�"�<�\BC��%���\�_���!�i����f1���v�R	-�h�I���(&�/�9|$�_���һ���E��;N%e5�<�m�q'���r��d}�[*���R�k�A	�x�&3��G�����8�iθ�S�bY�y!+iwS^�:��1�Q��#it�4�#���}|���4��h,%M��m{<��r�ML-��V0��dn����x��>�t�0��d�^��r�B-�����@7�\�S�<�����X6P4y���r�omՔ�($�PP�R` ��{]�������BvW_�_���x��=s���������}�VZ B�"K�$5j�Jjs%�4Wl~���j�W�%��:}C���Р�al���%x��ܢ���,�*�Z�C�����S���X
�0Ps����XJV�R\&ԧ���yś�5�Х8�ۖ�4��;𻐝��~��>D�"Y�a�wM~�����,�c^<0�x�E(������Q'vnl��HPP)Z)AU����9ڰ*�������H�J�Np����.���bSH�6�nrncL��{��b��j�	��3R�/P�����b-R��ֵ��P�[w���O�f���Y�C��]#` ��!�P�i��S_�Jኁ�d���b
Dc��\�ByP
��Ϩ�c5W�^���x����" 6��(-iC���V&9�O�qk��.�W�l�x�[RECљ�����.+�ٳ�2�0�����n�[3�b	L����d�sl��G>8�
��Z~��~zxrO&6�+_�*j��Y����?�U ە_j�gV*�~�u�X��Ov�Z���KD�r/���",O(����啳����([�ϩ�wM��@���[Gǚ�7� RW��R��-�έyC��-��;�H����F�L����G� ?�
g�!k2'��]�J�|+Ф�Y��Z��'�aJ��[���,�d��j���	��-o��fv�}�T]�V=u/i���]Q��'��]Җ���g|��B*^�n��V�e�~�N�S���'��C����
�r~���.&�Ra_txϙ���7��ri*!GZ-=�e�^$��6�ӄ���r�J�SQW�.����z<o�7
���jxJ"���7����=w�j����`l,���|���p�O 3�H��'k"�tڮs�s5��F��=Pl�[
!�
���M�&��OiJ��?	\ŷat��Ul��c�UU��/聠��N��Ӣ�-��)�U����g��}��rYN��:�>[����}��g����T�hh~�MFؔ�;����_�y�D���@B5$�Z����jDkU@��Dm5�ɘ=t�<ذ��)��v�VЖP�Ñ�+��t/zi�`)_�b��q���O��r2��z��r��"Gk����bt�¢ ���Lv��8��-�-�k��I]I`�z4Ba}u���K����'��r�VP8xz��¿�M�'�	d�?�S���NWpi��|��Nl���V�:T���6sn���2"X��PB1	:��� :#��۷8tO0�����(u�췩�p�iH��p�5\G�u�Q6��� ����+̧>VW�� E@ /����n�<��FP�����cč���������*xJ#M"|�I�<�R��,Փ��_��FF��{t��$Չ���vI�Ӌ���o�C��E�i&�	_��m��5���
���OD�O��A""�H� t>w���`6s�����N��|"�<_�|O���T2�b���w�$T ��_h�B\5("Q���&�Y}��(�.��Q��"1&�7��$��1M�*%��A�����)���&�U��R+��jM^�]���DEL��ԲU�)�IW���p*l	�v�N���9�!Q9EJ5�?R��fp�4���P��;�'7:*�y���?���(S��L�t=��3@�9�	�9��o�h��T�\�M|�E� �4P�D��Ҧ3��|�
E��@-­�����������jS��yD����������;H4#��>ž��L'��)�j�2dM����7Żyi���������3��I3�QdQ��-'6m�O���#��.���fm�%/���֫�j�p9*�ɇ���ȩڿ�hO�VAG|{r���a��s��gJ���E���$NN��<y�!�d�֗Rp�&F����H.�6�}kS�v��殒Mrn����5-;3�����@u!~~k濱y��T�?� YZ������5���a�'l�:��u����'.aC�8�0���Z�ӻ��QקO^�\%�;�+�׫>��0z]n���f��ر��|ǶRs�� ���;�F�^5H�۟�7�tl&$��w�?>Q0�:�8��AQ�����'T�� ��P�Ov�	�;C��z��O9�K6�s �z�=�d�j���L������7$��XVɣ�6Cܤ���{�c������3����UՏ�-Q`muY Z�C�m�I�
t}S�[��
�6>VN4�����o8K[Dݰ�U�)�F[A\�B�h�+?�ͭgk���/mB���S��W�C�- �zEO)�i���]���W��\�|��j�"�)��:~�.}((��}{0՜�X��)�$��:Fi�~��P��t�B�����p����7�)$����Ƭ�tE�ѱ�T���e(�U�q�&q��0�����D��`��o�R�$|9�PUݴ���E��������#�J�簈���-����	�*?/5B��ra����sq��bqǏ�H�ޭ��(���T���J��F���]�P#a�ձ4	���ܑ�����`Jӆ"Mcf��l��]� �>�cq@��oy��k�ҙ����/Q�(oEmϖFk�`@�� �f�&���.�ߨ,p��{ED�M����N��F���i��i��V�;�����o�_(�@4+l�%D��'+���&?Afg�3|�:�b`�j�`x����.������I"�3�x"-��+�� 7 y���9�B#I��R��K�>D���vi ��䴐�~�3ƫ��@�s�(��S�u>�rK�I.���,������T�טFL�'����x8Bu�-Y�j���/�N���l���� :9|j,U��b����eRX#XD���!=�۝�qR��SI	�7~'^�Z/�w�@�@�͠H�����5�a�,�>��q*��#�bj.��W�瞯[�l�Ɋr�K���g�	g{<מ,��sW�QGB|�o�����OD�ޕY�:�,�Q�
���Jmu��hDS��@`��E��_�0��Ԙq��v���n)FA���E�2$�.�ɩ�Z��Eh9��͵Kj�Br�߶W%������	�n��<�ƶ����K��`���������;�M3�"����*}�U�3�����69<��Ճ����廯���U�|/*��7tPVI�"W46@��������<�1B�q4U᠟�π	M�u~#���9�F�/=�&,{�зE��,��m6\����CL �K�u��0���"�T��lF�QTx��g�ۨ������:Hk�����͋Ω���@��R�IG�uZ��\�	~�l�Wk�pvZ��эN���$x!�$���eh�r�����*�k\�R�(Y8���V��p�+ϝ�:6��?ǯ�\iA�}�Af��X/J�d9g����p�-]>�곝����2�N�)̤��T>F�I����H�!d���s����~��֜� ��+�Kk��I��{����H86	!@�0�i�x��Gqm��u�dꎀQ[[��o�ө{���N��X��<�R��/,�D��vU��}U�N6n⫆��C��s`1�uo̧� ��:�v�R��;_ټy���ǎ��Z��EUb��a���1{+��>[�j�̇J1^��{��b�	��������D��>�<���[@�)0 �N�u��+;s��<Y.����i�7|�%�����2u{��S���kCRt~'����=@��uS��F�1*��>_jW�i��r�������'Mp���S�Pv�ѽ��/�4V�ׅM㱈��d�B���'����8l]��N+=t��W�w��Rr��r�YD.#��&Gc�9��8c'��t�n����,��æ?��Y�'G���4v�]w���l�b&i�=�n����k܍�ʷz�A��[����=T*А.�۞��j�e�尐��_����'�ұ~��o'�{� 1CC�I$�6��Ϩ���ao��*��Y<�i��l�ڱ;��=!�UI���:�[V�zO�;��"<<y�?���U.V��?=�u�)3�nEJ(yD���wSB�׮(M[�]�B����x�R@$�}�����aQ���T�B�)
Y+�8����ؑ؁��{u#��H�T4	�vp�1P�7 h����n`�:m\_�T��Q+�~����������I�Cr�su'��T�U'����!2Z@	0o�X ��5����`�w;���î␤ 7�^�I��s��]<�<��c�	�K��/�S���N�F���q�[���A$�� | �U^;�L��'�:��KTk��g�2y�ǿi/n���KZ�;	�h����蘽 �ߦL.��}S��ܺ_ϗc�� �]7r���>������h��C��m�2)�8���1�H5���v�޸=^���v���q���ə��/��s����n���K�B(8���}ȭO��L��B�h�V]fL�>��C@�0 �m�aL����X���2BNV�;�L|~�S�5�rჁ������Q�x�JcTCk����]JNrB��F�K��jҹ�GmP�lܫ�~�g�% ,�lhcYE���� *���m.`�pG�q6TXC`��$E�M��feU�a���_^}�"s1��ɧ&��D�b�g���f�U����'J��1�80pR�	��<G�܅������?a�VO@Uxd���E�S���ĵ�^��Xe�1�I3 �>8��$�%�|���[_.]S����	b��Y��𯯛�5�ZG���%)�.��za�� �_�,ς^���+����J���~h�/_RhXسC�5�� �[�i�zȸ�K\�%��T�˶QCZ�o,Q���3�J��L�\MA�_n�^aU������NAN��) �אz�a��q�Ka���ċ��3}��'ޖ �6(�yB+��k#%U���U��o�:��K�]����� '+ML����pbf�B��ܽv��hZ�g�� ���0 ��'��&}��|�l��
@(���Da8(��e��o�\�4z�R�_�ٔ#3�MJ�<��L|ڞ���J��#�1��t �<�����G�O��Y� s+���əx�k�F^������r_W�W�m��zc-�F�qBO�=~uZ@�)J��+G�u�] M����-ye�������2_�U�]�Ū�;h� �/���l� A�h�N��^<IF����t�x�eE^�H�l����Y�����(�s��J��F;�n|�D��K$�)үZ����� ������{���{bXLrN�jԖxh�LG���P-����Q����o+�dGt������e�$��$}��Jc�[Gx�0�%W���K�᬴醂1�#�0�.���ܘC���*
ՕQ#��'tY�yd�*tnz�iӑY���m��<
�:m�~�Bӗy�J����C�K%'Z��7~\�ރ��2j��v� /���$��Ū�$�F��ƌ?v���uP�!���J(	! =����2�on����|��ۅ���T�q;V/��r�<�%���\�)�q���"mi=@"��Χ����ꦙ�KX����92��)	��g��~*@�*�XSItX�((�%d�01<ܡb�;L9y-B	�x	�Y+�(|@d�h�p���{��C�"�M:G�ŗ>�C���������w���9`� �V}��r8X�Mu�S���g�ً90��\�;����k��8�p�x�<7�1u6�b����sQF.O���fMKQ�Yc99�hh�<9�2)^~�: ���1�M�����wց\�'�RfJ��Ot��޼x3�qE�%"��Ah��]����O}��`3/J4����=�w�D��������Oj�+I�(�����b��O�)"��+��idW,g��v���3�F��xd�,c����-6Rw��t�:o��� ���Pļk��YsD�{�Aq!O`x4����>�'����/�ud>�3�03]�R�x��]w�Q�����
��\��]��]Q������X��Bn0�
׍؆j�1ݯ�|ԏ�wPl�Gs�Q��6q�L���U�܅�;��=/r�`�C'a����;�\�s\�v=L�qv��d�y[dy��+;-�0�<�<�"��oU�K_k_�l�~q͹셐C+HV��!�ڢE�-$/Z
cD�mY��ۆO2�`e�p�1|����u�
���v�_�8?�~�8�y����<�k�z	�@�{E�nt��K�����=Q�P@@��n㮙a�H�3 '@���3�+�Ň���wak: L�����
6��OE������d�o'I�	�R���?�7Kߑ]
����h��L`�wI�~�p�5�����(��zd�������Z��
�nq���%�5c���\�c���f�A�
Lܯ���`[�f��K��u�Km۩D�/AN�&�D�WTsv��'C�/<
�ҳ$h�P�5R!�В]$�5A��6j�X����K�E �?��S����hD����eH�#5�$�MC�xT��I%	������-�z,��:�a˳v�d��p�aB���m���ݏ|�Y�m���T,�|z�15i�f4��
����)&���P�=��;�1�N-����x�����.��BI�
kb }ʦ]Z�l����V��Y���Y^�(�o�t�~�N.�ɼv�u� �Vwj��H ��F��7�1
ڕnEW^���g�G؋��6�_8�?�_TXN�KUdA���Z�!	I�~�92u�̓�F(�VuB�Q���+ث�k/�уƓ�"��hr0J�����Ob> ��֓F7^����y	p�|�Ͻ.���1�T�J�^�R���ͫ��^����.>T�!��#�^��ϐJռ�`�)�IIa�ν�_����i�t��C�V�2�yB�g
a=����ȑ�q���"���d����u�~7�T���ONFWU�i4�`�F�%��)�s���{���jo|�%��Ey���aܔp�%eag�ҡ9�XՔ�ձ�ѿ���8������l�_��w�?�0�=¯/$��"�ן᛽m�[X@��η-LY�MhU�'#:��Y!:��D�%���}c�'��η}���؏ϥP8�ړ��`S��P�(:��1A�@����[]Q!{uD2�V;d/�|�.ɝ�꾐B��[�Zڡ+�2_����2u��i�V������0��~�5�*�^-!Ȕ9&���(*�����k�O�FT�&�>7�i�s��
��K� ��$������3 Oݗno�$����2��%ojD/:�ї�ߐ���?8�Y�(�X@A�jT��0�9�6�
��Ƚ�q�����J~���@Ѳ�ԥ/��c������*!^� z���eaJE[�����(�t���RLk���ZZK�)`�͞i����2���\��k���F���C�AD���D�#%�S/�1x����݄�&�g�SR��S��"/e��~���@e������1�{��N��.<���ѥO��ԇ��_��~72�ָ�A��%
�<8[*Vr��v⤚s����K):�ѣXԝ��dI�x%��m�ܦ�|G���(+�Նe�-3ss�\^�7���%P`������1�\��z�� �#�im�' ���g��Jmlo��Kz/ީ����	�HM��H$D���[��]��&y:s�!�k�՚@bָ*Eh-f�M����!��4�jd���������X�kG6�L�����z*]+��#\�{HnJ�۰�w���2�TKr����3���ԕC|R�G�޾����j�{��(7Y¡t�Q��F����Ǝ�}]Z�JV��P�i�u��TrQ�(�Hh�D{����EI�B~hʻ��G�d%�d1�ܶ�{�i�wb�ߝT��-a]�2D��<��h0������kޕʹ�M���J��*�9����N�<ٽ�3���m��)5�}�]��ˬe���F}�U��Ha���{{���/���{�(ۆt�K3���<(�in��#����-��v�I�8�(}ar��iωt��x- Xʲ��ō��ه�8
�x�,���������h %{�tD�[V'��Ѱ.��G��G�-��'X|]Ť�S�������v�[-�Xf�Ћc����(�n��=��ܯ���F.������[q�r����������W|>��
�	�&�#���B�����M�"���ΒX:��&ц�,�]�+��s �����	tR�&���Xq���̬�|^1%�
L���<Jl��*��!4���
>�)����<|�Kh27Lܡ4�����;E���h����� �b��s4����AA�Q���WU(���{�p;��M;���||�
�a��iЄ[V��m�^��\®���ӳi��n���4�'a(4�eU�9�T�
L_!(���Np1(�¬}@�iDR�0�X���c�!P��0"}=�!��۞pA����09��*��A�������ֹ}������40�����k��NFa�O_X����l<��������d�/{h�<|� ��?�G]4J,
�G��[D+ڴ�C�:ԯ5�|P���]�]�t�S�#5��-����O�T�}�Ր��[������а{W��td��V���\�x��@�X��.���,�Dv�:�V<�8(��>N�P��o��^Sɔ����uX���k1D2�cV�3`���Q��yb\��4��[�x�uow��Յ*��i�ǂ�	��*�|��)���g��_
���C�(?�?aa��Mʟ f�&�Q�����_�(i�FD�"�q�=�	{���oe�+��v��Ì���ÄfI������xjt��v6�޷�Ӝ�����Y����ObJS�e�[���['��z�p����ы,_��~����Q��Ƃ"�4(��m\��Q�>?)�$���b��Hi�/7���d�<sW1Đ��R*�� MBo;�f�I�Ø���j�S��VH�����;�-S#�X�Є�� �(�І(�M�m�w�Xh�FT�����ER�]T������L���b��&�����o9�خ"� N$��[��t���_����$&��[N�0��a>H0W2;��Z�lJ�_m�f����i4ܿRT���ϵ�k��&W,Q�!����{���`Gӝ��ʬ{��,��I=|�[�����K݄��fO���>W����v��pܰ�2����}�6I��dX��dK'#�VtکJ�)f�0��A���ݣ|�|b�8��( ��������*	������q���[{�!����j�	�l�łr���E��o���b���v�m3]6�X9���]�9\+&
�Z?�	���8���V/}�=��/�\蚢T�֌4���wmGe�+׿��oj��YB}v�I�sl�����?�!B7ać1�3���g�M��6��z��fMj��G�Y��>XY�~��;YpT��J���;��w������̝��i噴"֣�R�JJ��%6�LD�� �~�$c5� �un���D�ȷ�n��_�Y<�9�8Ǐ�t�Ӿ)��P.]�t��e��~أ^�i>��5���kl�_�_��,�t-�'��J�}R2O�zBQ���=3r+��'��!b�K������\��瞸h�r����.^��ȽzF"�N�`��tY���<�>/�M� !��AԐɉ�@V�����V�������l]��)e��/B�d'��Ȁ�,~Yn�L.���]�{��U�U�o��d���aL�FR�<ܣc����z	����N��5Y��\`�»d�𰖼��\��I\�P� ���䞞���EG|�G{T	O��x�~���e��������H(w�&E�^�׈���t������E��GW�j9�C��?M�5пĶ����=Qd�|$v�/v9�m�S�9~^"��/����7��|&k���z84�y�N&����Nax��v�J�KI죇�8}�W����Br����@w��'�(���!����E;Y:.�9�D8!��A�;��m���L�X�C��?ʮ��6׀�I��0����*���D^���$�y+��3��K&�c�o�#�?�&|-�r�g!-�e��GN�%{.���LV�MYc�#� =�9X���Ys�KǍ1�'��/��a*��Vك����m�9�N�Ys��L�'�|�q�x��/ȁ�;���?Z��5�l3�V��WV-Sr���1�[8��i�WF���k=c�g"��w'�nZ�i�E��p�,7T�'�����ܰ?v��]�m���H��Z�٣F�2�`9����|�AR�����)�Z�UY�u������<8=� ���?�kփ�` �S����3�0`��j
t-�a�@Q��=Z0����tRƗ��̗��p����ĭ�[8o��O\��]2��Q��$���z��a������#B�%>�)�.�y��O��).<�a�+��V%�W���P�}�K�[��q�����$��T�L�/^w�o���`�7������l6ڡ���)�����@6ʨ$tq��p�/C�t�r�k�U-�:��VYl��5W-��G����4�M� �C�� �8�[v%J-N\T�\�M_g���~�'��E`������~�4��vs*�u{5��d\������ 0�.�
��̶1�����l���"Du���ؠ�%ݝ����^��1�T�8A�U���,�몮�k�"���������l[d9�>��źq�U+ \9�+�gma4��4�M��/�ʲܲ궱������N'�Hû��V�ۈ����l�ѡ3Y#���B�jN�9n�}��MN����AZ��J���(}@G�����Ǽq����|��5f�	VW�U#�1C�Ɠ�^^S���>*��z�&u��yޱ@ѩ����]���-@�p�<�D���(��fl'
���5�o�}�[+�	��-!,�����׌@�ɔ��̮^�"}��O���OE�Vs�۷��K��E���B���k���t�<�%`R�5����|:[�s؇�2Xѣ�o�j��궟�Y0�9W=h���Pp�jm���MF��V!�o���Jp�D���rK=��_�+���Q�uz/L���܉�i�S���nݧh�}�Id�:�|�=V�s��ԵF;��c��
�.�J�R���O��Sw�]��r���s��
[i$��2<p��(TU���ho��g��"r�%����ޞ�������Hbl�n��5h�|�����<&���ˢ9������hc�����ѓ��R5�������sچ,-��./U�л
)JR���y�F�x$! 1`�;������(���]?��D5�^�E!�ۢ�ɢ r����!ZO�z�(9�d���9���د�غ��Ә0�����FZ �IG;�B� �A3�\�