��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� j^ꘜI��e�cA�ҏs��U�eM�{E��^���4NqM���(d���˙�Q��������"������,�Ŋ�+ɺ#��}ϼ�Ez\,��
r��*�x�̱��N��TfI�PO)J�N�i�C�+�C;_�PC��,�P�On��E��;7_�d�j� �]�a�c��4�c�j�X�� �8�N�2K����
���_�g"c�l7�M��2FWa��%�{�H*��CR���b,�evmҬ:�҇���0�Z� ��>���w�M�*��jA���U�H�0����U�_~��Rz�mѳz� P�����oAş}�Z�|9m`�~#ť|PV��9������!M �7X?z�8M��'��t��rǹ)�˨0��a&A�\:�d�F��݃�zFMd],G����[l�kA/�<?͠����`���aS�|E���]��'DT�1!��DJ�'�Eh�O&2���٢yVuA
 p7�^ar����>^z0��5�ZC-��c��
C��
��4��W���vJ{�Juv�mjZ+���`�d���m�H�������r?n�5�^��ʡ�6�����5s�����j�ߋ<	R"Fi�):���ë  ��M����o�������`��D�5���7��s	ɿq��w��[y?��'b'���<t�vZ��/��7�c�/�&~(��F�K2���MB��&J�*�hO"8nI>|��E2����]����AQ�)W��\�)	�g&�XΥ_YG���]Q��u?�ԃ�L	����4�9�
\�͕��j��8n�{[�|��1������J �����ر�zk�ՇED�
��zǒq�����SPc�!no��(>�ב{{`���hm�(�C������G��#5�O;�ocpD��H�7����L7�h��6�3-ݾqPi����⡹1m3Vox�T�`p�D������]�S�:��4t����%4	u�C�碏��b��g!��s��H��no�m��u.��͎�6 ���A��\@m1��Z(u���G�-e��m�7wC?�Bn$$�%@×�|�$�g�٦��z��U��X�v�Ǎ+�WG{��Պ�c�$����LC������]�LDT5�� �<�Ѩ�N����Qd�8��뛊=�x	��P`%�R2<���*��l?n�ݓ%y��7$A��躰�㲁s�7
�0�xF��<vk9��H�a��2��A&�m :�"u��S���{JҠ��rj�KsH�Ծ i�F��%_������)��f��}z�𾒘�휎8�t�-���9�� &�e�$�I=�Je}(ԛ����z���V����I�]����h�w�zw�y�A��>�?��bK+CV�n� h�.2޺(YT	\A�|����l�y��(
��G�g�.�;���c:s_�jR�����h�*����-�{�D��-ʦ}��2�^=.�Pv/ji�$�n���.��@-�����,����%b��Y��G`Я
�HM��.�
9�'Z?����f�0������ 
���������RĊ���� ���l׍0�=NwR�OĄw�> @��z]�8��|C���GCId�܎'�a����e2l���^��U]D��X<HtX�ّ�E�E�<�;!_2@�H4����y� �U���nX�\���G2�B�<�'�0�����%dT���g�4�ֱGj�^O�U������byª%K5x�Ն�4xj��,v� �C�i�9�aA���i���LlJQ��r�uU`W�-̱x�g�m�LkaP��n�P!yQ�5z�viU�`�O7�G�ݛ�Syw�q
YߊL���JG�k��
-m��Eɜ��(��*�)������T�0�6<���R�*?A��	{��p�!�U�O^���&E$�r�|[�3@U)���r��!���=��-/�P�N� w�NgZ�3�,*U����1Q��Փ�k%��fG}r��:I��:��ⶫޫ�-�'A,���"�N�����tc?;���n��u��ˋg96����$�pG)��4�p�4�ِ_a;�gyo��MHWz��������bn��3 P��Vg����o����Y>m!�0�_��	</�;�H�'�b=�`�<����[���?��Y�X�v�(���u���|���`D��D����non�R�m�cL� k?�Rb����6�~o���rm�l3T1���,b%���y�J�*�6����_��6� E������x |���z�p���V=$�svӋ難���T�4�������	�����|6���W�ù�X�c��N��[xM��)/�~��Z�����J9���4�W�gmw|ǒ���������� ��^�O�T�;У�K� ����#ڈ����]�cg@�S۩�H��/����i�dQ���<��;�.��!�]�K�)Ɯ�I�������Ż~Pp,.؂��)M�"�,�Y�ͯ�l���w��ߞ0�ڤ�ᇇ��h��� �������b���E�[�9��SGg^ngv�x�o����-���U�.t. �{��~��Ѵ�_8/��ap��E8��� hPc�k���] F��^��X$",RT����]�vR��h�'ZJ�M��26C�8��v�7�,F��*�8��oO� '%�B�*�#f �یm}*T�Q���9G�� ���1�Y-��9�P,48@b����Z|�X���0��Le�4SNT�$�8o)��μ7����Gz�H,9`�;�Zk/W��9�`�z��d�Ȗ�L9�1�j�_�Q�)X�p��x9��iy�:����ז�^��p��I�G�k�A|��ݙ,p����6L�3��#��%��7��h�ˬ�"|����[�5;�bB6���(c4&���(��v�`z��EzRX��ޫ��8K�.a/u(b����׫G�?���GҠ���ݎ��sdʭZ.y0\I��4�Q��0�`�[`�ϱ��
���k��w9F�z_�awf������6.W�̑;{�G���^�[�|�2���
;����.d��a�H��a��������!M懐xv����"�C(��Y�����F��k�6�Y��M���]�M��i��;�Cϐ�b>�yD��=-9"Š\V���7ˉ�\q����@w꽺��+����i
�ƥ����g�W�9�&���c�ո�#���L'�gv��%Z�Y�w�����K��!hӏ�f� �qtn5�D��i2h~ Ƥ�:���� �)+��-`��Sah�a��߀ڴ�}�
+�ܫm�~��	 K�(^˕�B:�b�{e�du5�
B�)^-^��D:5�4_w��y��1���*8{�_`^�>�p�s�����)@%
��w�w4zuB�o�?�������o�F]��xʵ������D*�s��B�t{?P���@��"j��I*b���*��ȏ�_7��$b�	�5m��R�t��(�o�o���������reK+����{C�m:Em�g���$��(K43nc���� �HV�_0���c����k��	{9��s�'���|��(��GH���= P iD�A�*���R`�����"�7��Vqx�Vb
���8P�|a��ʦ]NB�A��c��ؤ/�L����KKQuQ�}+�b��;��	��E�y\�S��p?�?G�5�Щ.R{J��+^.LGL�f���5zfP>!�*D�g"�r�	�N;Atpn(8C�Il����9�"������-d����+��fFܴ�INy��6��x@�;2�3
�����0������r���']sd<b���6�KjWu<��i��M�Y���y�8C�}ڧ�a���Ţ�S9~ �G�� EP@���ʶ�#D\�� ��t��u��`V��ZHp�5��8꣕��7օk:�h6��U흞�\W�W@�껚�'�4��`�Z�zQ,*��L4�ɵ���(�x`�ɣ��g�gT$qatp���vc��V�������Q�v�_i�0�ϳ����F�2�1_"LTIwG	��d�ud{���۝4�1������쾁a�$\Ӡ0�����=ޛ�N���q�4�KZu��[�	\��-�d8�n��ۤRIfR� �8��W�f�}=9[G[&��k��S�a�4�V�aG��AepWmg����SB�M�+z���Z*��y�`e�FA ���r���6�r���K4g��;������������ɡC�u����iRz�~7��e/�M�dN�4���o��@YRR�޴�����Seֵ��RՒ%���dl�n1�]/���1�r�h��fd�⥑7gU۲d)��	��1��y�e�3��ے,g�R?y�C줁��_�0Rw����N�kU�_�u��#��R	b�������Q��~x�Ȳ��_Uh]��O�m?�������"�fg𳓉��t���}��ƀ��mN�dݾ��	�����bY��e��ex�<P��e�="���q+4��t��0�P����)$�^y��f(�jD�q�:�'Eag�dS?�`m�o�S�|�>����^,ٜPr'�NiWɲ�u��+��4I�`A�/���^�ԫ4e�#�����\���>�jt�C�
��nB���C��[���Tf �X�J9������A�j�EZ�����~��^]&�v�V�1d��*>%0��sA�\(����gT'�{��}����!+�þq��`�E�9Uv�^��eV��Z�!�qi.U}�1��
q;���w-�x@����3��z��J���J��yb��B9�:�<`2�) ��P9����v����x�v�H
�GO���*�*,��2Db̰������I���-G�#o�!z�� EˮC�巺#Wk;O+���:O?N�>�N�c/�	�t'��e#�=~W�傜�,q�r~�pf��l�Y�
z��KcP�����q�?$ �]@MO"�d�R���(lE�d�S ���*�ha��ޔl�l��貈6��a���T��o7����y�)A�ߨ�",r)��1�H�-�(M��3��f�[�����/!�?�[���a7܃O��j���U�).��a�TܗY�p��`~f���0l�K)εtA\�iPnD�7VτU��zȊ:u�h�_�N}���b���;���pB8�u݁EjT��x���y��_��z����U����0.�͉�fi�Gv��a�9
9�_�(d\L�:�E����3��%�����M�x�.��C��X��J�*i���ܽ�����At��*��OE1��B�2o:_�����ј���c�����Q��Z�����,55,�!�pP����p@�
_�tf��蛴��ݲ�E�{��x�uv��`�
m�48��)ٝi�E�%���z��+�N-�0��!�:0�=�7�;��gǈ�Q�Z�B�q���q�����?d�Ip�A��b��m=쾃L�Y�9:��1�|v�؎�5A��?A�!oQ��|�KJ�UCd7�N��.Q�ҩlkA�����ʨ{}"�_��Ф�)�" �g+���t��J2Z����7�������4�~�7���&5�h�1iu�*��?�����_�ūp�X�Ewԏ4�%/L���*���F:F�+4�ոq��⼔�r�=�e����D��@ )�:.�D���!���B�����'��l2���Qw�Z�a��X���A8����_���̒;
`������4�7~�~t%T0��[qՌ��D�����x������L�Ƕ���U�(�_?L;�ֈ�$�3P�m��GF=��L(\�������߸�a#�R���.�gv,�"����Z���.�^;�:o4)�>Di��#��Akg�s�N�n��/�z��6�EoW�ek�y��G)�J��)Л�SmL���7��w�f{� 8Xx�U��舨-��-J埚Kނ��d��#�Ξ^���K��|��2���ð�m������T�������u�$��+B���d$3������!%�yt�^Ak`XlA��:1��U�
0T�KɄ��B�)0�-�� ���hY�[M��(]�j�2D�l�B�ۻ�"�Z���G�Aӽ��x1�'dQ9�e?����	z���xAF^1#����2<Zԍ��R�O��?�#eMk�[2����6���-��c��Y�b�L=��{�� ���dX�Ar}��ޛ�
@��[�&�*�,y�`�G�w��FՔ���B��e������Ƞ��.��A�q9F[['1ݐ
��\|����t���*}LW�����hs���	�g0I�`�����{�G�o�@c=���}�;9@o�?����Ki	<�y�/L:�v�MG��2몢"s�
�y�6�d(!�ɰ��u��:gA�*Gi��C����p;,����X�ގqD�f����-g���_|UP�M�A�;_��\���,0�e,�펐�bN=^�c����y䲃�l`;{-�ӝ�q�eso���紞zͱ�^Cnÿ���Li2�����l$��g=��D���l��S�ЯC���r� ��؅D���"�ެc
���Rnd}���1Gr�D߷U������d]a����9���>�$&�⿪.���$�>��lIr�WE9zV=�^���������uoh���Fzߕ�;��Ŝ֮{��>��S����������Z�ZqPxw�S��t$��0]�m�F���+�;�؛u��~��4���Lg�W�=�؎P��|m�{��,�����I'��#�X�2 b�Dev����p��+���Um�tlZ�����N:�U���;,��=`%�A9�����-�)�[x�qyI��j��������{q��r��A��y$p��W�|�Ӱ��m�v~��`��������<>�
�M���5� �m�4��_�f,\AU��9��G��]���L\�����W��AA�DM��d���ZAN�9�)�%�b��]t�6�mx���r�TXUΝpP0�B܍'�a���'�D[eAbʂ��3 wӒ0O��}��7�[K�ol��^�g�#[��ۑ��T��\��&DH�o1�{	Ww
+A�����n�@L���h�xq6�O�l��h�rT���On@lPz�U��H��w;P�k7�tr����o\$^ҙ8��P�	��'��@22i��md[����G⋝t1��F�b0!�k���=�CA���X�W�&��߻)�1�]d1yM�r���z|�+
rD{��)�<Pt�؟�� �=T���X�K;�;�Lv:P�%3�,E' �E5�z��]aZ�w�I4���/��j��0QJh^�c�����ү���0�d2�8�Ƕ�:���hm,�	v�/�..�1g�]\F�};az�|qw#����s�Q�G��~w���[�wa�V^X����k����|:��3�Lp�z����x�fo���B9�7�Z�߮�^C��.fe��m"��-S�J!.ב_.��[DO��r����ݤR�}]���Z���#�L�L)����������~kbP�vy�W��"(H�a���jðO:�pT�r��]�����ч�e능W�*Ǥ0e�,��� wb�UZE����;����3�K�6_ZJ���U{xK�2
/��8i�=��
�;&(0�v�q�~��V����`)�vYu�w���]��D���cE��Fږ�����ʬ�J9�������Jc���
�,���&���ۦߚ$q��i"q��7���ܩ~?n))k�r����:���z�h		��3B��_�G$%���ގt�>�Y�E�['��⮑�ͻ�����Ǔ��MQ���S,��`Z2ɪ<�ng�d�[[Բ��5��<���b�5�@`�����x׬�AI��yٔ���F�/�-7��YN;�tp�n?olz�@Ց�0���@�:���{N��	t3p,�F|sB�]ʳ���A��]���e+�d��c߃h6��|_�<t����
~�{�9!Y�4ר�)AV�ig&k���k�g��d�H�x��tQ�$�:h�~��"|��^��}_��! �C��LYL�"�΁D�Npi�,2O0O�!�r*�Pu�G��P�C�[᭷�P����(��E�=�6ap�+�_�0+*L��_�rF����A��gu'���Y��;}N72��з��e[�Ն{��}#�7��`���	����=�5G�'W���Z̩�`��M{AmK\e���䟆���^@,#�W���8%�N�Ӳ�@���7�n��Q���U�V�ܚ�k�">�P,�MWR��Q6g*����v�$�8S@��~�*BnM������.o�Y�0ؙ��i�#ݨ�VI��2čs��M�ț��jn�&_�&�x�H�:�x0�B�a�E��pp�<��5*:���]���x�N�f ���Yԙ��+IK�>4ZY�t��
p���H��BI_g��oo�*ɴx��Ý�Z|��8�*�8�A�g|�V��Ɯg�wR��;�</�sR�&txi�B2�ܛ�{~��)߰P���k!&\t��Q�������� ��(�g��~$������=�q����;��+j�Ї���w���χ���������]� �Ia�L�)�+%��_����òj���rHf^+:�Cӎ�c$�Raj�	B�ܦ��Е~����0)ƛ��HhS[P��,B��.|��JF����_;�^�d�wo��,SA?Oȿ�C��z��$D@�u8�HL��ٴZ��{~]K
k��U.�܉����Ѽtc��	P[mtHp�N`�-Y( ���WO!O��z�m��/�?/#bU�Qx�3#��ͨ�'f���\���D�*n�����Agh��DH;s2��X�WZ�x����I���P��Z�m*����	�D��Pg"����,�5�+��� i���Ʒ�j'v�k"�R�q˰We{�fF0ny]��SZ�^2��A_����]O|zZ�T�ՙ�q���X��]'��Mg,,ݛ���9"��ن>�҂�B�:�V3U�������D`y���T��?�8 ��}���=|�bl�2�bY
�.�xɾ�r��!����*��t�!��ZA"$�����|�n�էn�B�U��%�}_0Z���K&G���fV��PR�8]'��5⭥�B�����z�����K&ګ> �3�BF-3�oq^j'��숨�[@J��J�v�ۅNJ��G��b� Ա�]Kk6���Dd�;)��ΪŮ�)��.�K�^���f��=Y٬�]��'�_�����{�y0�ÿ�Z0̪�Z�7m�����\�@b_�4p��UQ�G�ӚL���`tq�\��"N-��z���)��PVj�6OC2j@�?�)$�����+�6��/#G�����F�<0�l���~�'��K�Ay<�Г;��`W�]U�oyI{��i��m����f8KƞX�[��.z����oA>��-�ӹ�$�# \�Xf��:C6r����5��X$~���&+a��vC��gW-�r-/�9oe�>��m*�x5����L��5s�%�6ۂ�@pQq��fT}���ǥ�,�
�#/��l��`��~۷��USv�6��~��H6TۡD�6	�!���B0?gM���8�{�b+*ǋ���
�{7��N�d�Qt��� h �ǚ�jt��ҭ���37=����6����f�P	Is���_�|��E����LvR�@�P�0���/�<=HQ��]i��
�01�%y�w��;�>Vl�������:^��	�?�۞���h[�/��ij;�=={�2W��֠v���ˣ�#��]��)ȗ�������%Y��+�S{���R�q��b�z����Kǲ#X�I��p�\q�AlU@���5�Y�S�}��-Q,=ee.�l��&�C��p�$�g=���gLݗ0��F�|��FIaR�A�Z���\Nɜ�Ǎ�����Bѵ�^��NiO��SC���b9Vl�HS̍�Ig�_KY+�A��١vtvҤ�����`�(N^:Ӹ��h�+�]��j��H��]?s띗��_r`G�����3e����p�+�ŀ�<A������Zqۡ���I6yd�)/��w�)�@�6Հ�� T��6=���!F��ƷT�T��L�����E� ��ܚl�gx�6����w�I�ʂr�Q���k�Ǒ�R+ �����t��bRɀ`xº@�����H��NIQr���X���ʔ���5�"�X��7�e�j�(�[�9�-0"�;�-��@"�f�SR/:�;o�+�̗�L�4�@�D��ˮ�.��L:��Z��Σ����6�����tC���KE	��#��0�=�ԟA��-��u�F9K�g>�_e��v�<\��A�os�}�W9��ev�.sE��g����%o�ҳt�cvJ̪Bc����˩����Y��	�`#:=ަ��0���k�*K��n>��*�- T�9�l3�4�Z���J����Z��~�e�a�n^J?���K��`h�6��Z���O�K�-�W���5_p��u�,�Jtv�-Q�<����$�tE�v�^^�؁}y#c����'�(��F�=��<���=�P��ƞ����˶�qnJ
������XgyF�O�Q�&¯��^��|4�	�|������0U �P7���:��V=I��+���5b̖�6�c3$u��	�������4W�h�;���HV��X�7sˇz8i[�ck��;�,C�me��c� �0evf%\�#*Od�P��O��U,ePGk��%9`�{��Lg8���7c����h�v	�vI{���ƽ_,�G==��8�^�jm쏧�6~�o���dCw�3�B;�d�n����%A�,D��tD�r���Imne�#頋���kO����s�y�x��7|�K�2 �;�'{�4t�OO���F7wi-ĐѴ'|��~��"����,��3lE��� ��oyYM��LU�j��H���VW�����[��g�xz��C��"����3���Ķ�e��H�t�IL�O,�Fk�vp�«�V
�춀����'�Ԍ�������<k;f����S 'چZ�Fa�o�K��+4L5iK_%�������:��l��P�*Se1A��%̠
���+sj w�5l��e{��$Z� P>ۆZ�}Z�V-9HH�2*:o��ۅ�D·�5��RHzq�uQ3(M���У���Y��x0~�|��=��G:�ЋnO5��:��$�~K���r���2��P~9
��Y�T6@U`��h0:�����`�!��F0xApw� ?���-����0��!�U�=���o�U!r�mAY�����HR)�_�g�(�Ƥ��F``?�)2�΂�5�zk	g�eٙ�D������F"58���Q}�#����ٱ�!�Q�,��U���k���چ�d?Wu{Nt��Q�l={vţM�@L��dxt��qp�n���$��g� �9�L\,��&D>�971�$iq�-�~!}Z���]Ӿ���$�5����[m�qz9�>�����w�`F���A��(Ϩ0�F5	���B��e8������vH~:�_�{,��7��+iܒd�9�uUg���<F�㔴tp���1��q������Q��e�q����f1�ί�޻�J�F���P���9�߾A�:֡�<��a�@߄N�ܡ�,9�"l�tR���N�wL	GKU�h�Wn�r��g��fe���T�]�������l"��`�E:�G(��b�{��� �["l~�J�Q�%e�@ ��O���rbv�FcI�Lb�G��h�(oC��>N�l;(Pv�t&ʞ�IbJa}�L�����?%�b H'L�DA�U}�e��?�m+��r�m�� 2��X�ׁ��ߏ�1�4�)��Y��ʿޓ��NZ ��N�Q :�)�2��P�Vl�XV՗%S-!"6
�T���)\�7����xE�F����W@�t�?�	��9vm4��>w q~|qK�Ɖ?�:K�6�>�I��%>&���ǜ��7A�}y�I��iNdy1�c�zhC��`�����:�8�
�#TϞ�?nU�/`�nX��^|�;X����x������]�]Z�:Q��Z?E]�
��ih�W��ygb>�Ӧ}��=�KN�l��qic}1���O�ӺL�RK��
p���;�S����4�%W�P���D��	2�y3N̛u#�lڟ�������a ��0>D�V�hTj��x�a�ub��B��s�|�i=�����Q@)ѿp���`�����A���^���[��u�^���6�ҳ��T05�|�8�t[�x\�Y�*���r�"��1/�. ���Ѫ�:�Ynɟh덬�����Z�B�#�x�!��jG܍u��ok$��G�,�x1Q�kWa,!C�\���1��Pwmg���ϻD@6��Y =�!Wpcq�q�=韡i��D7!4�7��8��Ν����eI�_nʿ���<�~9!��_[w=�9�b�X�-D�O����5�Y*���ZP���jS@�}[hr	��L~5�d"��E�Mvi���:xhh��g!��^����&�y��gL�ޒ����[ߣ�g��2�Ye�����R�}O�|��Uȯ:�JN��f(w��ؑe�3�~�l��$��-:�m�!�-�xi�!>H3,��; �T4���d-���_/A�p�4;U:���Ww�I���	p�/_ɸ\X��\�+�z�]�������=^����F��߂0� 9K2K]<��%�ۺ��
�Vk�!�ćv&�%V=�[����Ӑ<�������Dt��9q:�Q�XDr-㍛�;
�Y��)�t�V��LEZ��e�~S�&��s�>il����䯴7M�B��l%0gQ���1m�#sn�!9�(q�o�,(#��;�[�a�U�C��;���&eH"��3�+��9��헒��o�~�����'Q7���F T�B� Oi���Z��s��������� ���=�Biu���:�F<�d/���t�@m� �Dx�j�zw#���ڨ�2��`d��X�߮��WA�
�]?#��t�56U��q=�b���raw�ڹ�j�j`}�����Mgio%M��L��Ⱥw�W�����������@�z�3{E� \�(�V����� .W?��byY��� ��sG:�(���h:�˙���5+��ζ�n:ҁ�����(�M��Z���ؗqH��ã�7C>�O1 �8��i��Q�	-�O�oL�����M8u�j�f��j8N��[�ʈ��3�ͳx�Ŷ���e²u��[@�S7�:�����5_ߞ�W�`^�h�� E�>�_+�ЂN��c�f�̑G@�x�,��+��������G"�XQ}�`��.ò��,��.��'�i�]��H!$Af�*��Z]�)]�fM1Ň&:���j��m����cr��!,�՞�$,�5w.&i���������A?LB�>Q׍p,J�g�(+As.c_:�֕�\	A���A7�q��4�ǉ�Ra�]��e�4� _��LVg>�>{(�v�r �^ȑ�����~��������<7������u:A��˷y�X�� ��5սi�n�����|��+�u"k��0$s����y��n��[�l�>ʳ�*`C��7�z�g�z˦?��m��wE���`��o43�]g>e�Z�����S�8����_2����d�ki�4(^]�482N���DRè�*�YdJ7Ex��ra��p�V��B\�y3��Be?�_��� ��Z�+HI��I�c�������z�~[�;���o�j'Ʊ����- ��y&�[�qK��么�xo.��2.oR�����:����"8�aq��������[9�qxѯ+9������l;�;E����~Ǹ#6Q�6��~��Q�餇]Z�PL~"�� ��D�iJA�~��>k��q�`	ٌZ�6.�D�=D�Z��ur�R��Ekv����OZXM���֨�L�qE��Ѿ��F��=��Գ�T�(�qʅ͓�U^�b�\��>��M#�Z�x���m�tP�Lo/���,cZh,��MHAPWb�a�R�o���%��59.qg�	��3*��_�ci�V�p0u|i�:<W&!�����o���C��F�3?uRw�XQ�m���@U�g�kB���	��7��U�L����`�)5��;�g���].g�&�m� {4;0�;�m��4���:����2a�!�]o�<2��J2��`�q�\J|��v�w$Z��x�[Sx�'��O�iӖ���Z�G�(�ŕ�D?��+|�<�����HK��YA��c}��(�L^GRk�Qlnr6kx���A��i-�/��P'l8��Ŝ�d�m�E�ȋ��li!��ЛY��꽨%n��eb�^��W6�������(��[^R�(cSZ�֢�λ{��=��`;-��hx2�@?UzR;�ʘߣ)4����~/��c����=�Z(�{��_ngﶽB�*����+(/?�ooz���>�QR��H���կ@"x ��O#/�<,&T�el���Q�y�/SW�7�-(,��[yA:�tU�)�x@���j�v�l(ϖ7��;{#�1�d�6Z'#�:���d�P����Ii�|�o�j��0�\��T]���o�2�
�\˜��5E��=d@�������>�0.�O�qPDN�
-�3�Ó��QttI�|�#;8C�+��S��DCC@�e-#? �7`��g>C�2pY��'z0�H8�#탎��wL�B��o���(�`�E�Ψ�#ɲh79�@j�5�-#@��.
�����=p$Z!�͢7m;���?߾:�1���er|\ݺ.�Hf�5:�6bW����-]'��l��?x2��:�ч/%���dT��%���Qj���N�=z�����lB%#�	4!Dø��h+8
|,-w׵L�����NBvnc6�QZV��d�y>e�����A����XJ#+9��Ii�?�N,3^t�ba�Qq��?��R���x9¡���� �s^[j�T�e%�1��2)@����Cz���dS*&�$���2V�HUvPpߞP�(�r ���V�zu�.��d�3�XsT���Y����`�Jx�Kqg���'��Pė�J1���D�!ʋH�(��'��ۨ#׷��w
j��@��D�T�4�	W]%��zCE?O*�<��Z)����;�G�{ hƼOx�P�z��3��t"���ȁ8��n��dTHP���r���n"�=�3Ȧ��