��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-�D/�z�����K���LvݤJ�y\_�6�~��.���qۼ�R2�XڴvX���g����3����T�cP?��gYk��}�^uJ����"y���L�W�w��qQj����f�0�ਧLfB��)��(�H���-�aκ�i��k��nyKɄ�g�XA/9X���aV�dV�"{��>~��F���4P��� '��E��<�A[܆���ו��5*�`w���1��1D�����Ǳ	-(L��I�H��8b�:�7l&���vM��5V��`G�]�,�#�A�_�h���8F�����FC��m�d��>Pp�5a�k�R�L	]�(�C� ��:/�L>���Y׍��m,&W�nוRq���mt�ZDJ�!�\�Q,K�
J��q����?}� �� �����[��.�9�=�w>�s�	��L759H�C��F|A���o�|���V#�j�}U�ֻz����]�q+�����h��ȵ�N�E��;=e�Cp�' :�x���Ө7u�Q\V$�$�� �td��d��oCg<S8�s;��h,�0��Þ%�*��rcR6<%@�ےQS(��� Q�L��������'�!D��њȬ�w�u\FI�N�.�4k{_�(� c!ӕ%�E�a�A�,�늁M�=e��(SLD��N��ϙ�Ή{R(�/��7�-М}_��~7�%���#��(�*B|�l��P4���y������G'��{#�ԓ%����n��7S��pVD�D{���:m��S.}[�m�\��~G���j�ʛ���c���)�1euڴ����Vc�c@��'�Z|�L���Af�PB<�&T��(��{*����˩ԋ�R,�������~�ק�T���Ig'�5���0���4>�izC����mz�JO�ls�ԥ0�/�`^&X�m�P�Hrs�����9V�ye �2)�{}|p-��=��G��ۋ�<<L�7uyO	�>dz+��Oh�h+o�