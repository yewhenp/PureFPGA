��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ� �t;l�ʡ(a���mhέ�g�����a���E�� ���V�j�d�T���`�k���#�6��A�\�F��p@ YA���F�����ǥ����������I6�YV<)�OdM���B45vYڇ�h/I��U�q�KV�rwo�\p~��c�9�_�>`,u���������9֛���[T@Q�e�-�����_����ϋ����� �'��?K}\ ��8z�����*��uA4�g;W�"�Φ7��T�h4�K�.���W�Y
H��7�Bn�`*�oɖ�Fs��Q�(,�E�i�-��Q���剎���A���R�GS�-*ޕg�Ssu�kH�Y)�:�g�����R�� Hez�D�[��[��O��{X$2�?eK�hU�~�ҹ;�c C�?p
:3��!��+�X�vǘ.� 	��O��={`�5>���u�ع	�swQ�s*��,��b�7�͢*I���}n��L�
�[W&=��D�D�U$��)&U���q�@>�e�M��}�^��\;O�ZxN��`��<�9C�,�l���yA��<]����z1��5L�K޴O��	H�6c�q���'�#̚^�J�*���4�5d̈́`9��r�
-@ѐ���� � �=!%OC#�kЮ��4f~`3l L?~yi:0!�iU'���LW���5N�K3^�vxf���C6M�x���ԑ$3��v����N�_bՐ!�H���}��� sF��6Ih��%;�&�7���Ǩt�k�'7�͓��'�&��(G*1��h�QK6�r���.Xۥ����'�A7Tvl�P��O�Q��\fN�ӓ�s�U耻�׆�_c��譂^2o�W����¹�5� ��:^���l4�2H���y1�ӲW�}D���]cM�\%h�����͛*��9E�ʿb>��s��X�~B�)6ͺS�u��L���<`�BǦ�ܭ�ũrH߰T�!޹�����j�|O���/��h�r���QF���,肵H���UB�gW~,�~� �'+�B������mq��X+�`ԓ$���J�(��:OL&k$Xx:Q	�Xl�su�@"�,V�����ic#R�q�4^��gv!��)��v���8�%�/�2����+� ))��f��������$��t0�#�t��. *�����x(Q�H51>@9@�?��ȫf4W����^�p ܟW�nf�i���]~ ŭ�P�ri/jm��x���O����Re5�uچ�K��ҕ�Bi309�O����d}i��)>d��3'�̍Q�+�ayE`�]�<�'���$�x�%�m�P�l��I��o�O}�� >�{��I��%�B��� �M-�7�+pN@�Xl
Fxz��cKy�
�UB����?�;��%:"�KJ̴��$��xy+ٳ�6�Ą�1��j�:�6��.J�R$�4C��~u���@�2�I���"uij����)>5ql�A�J\DU#P�#�`�L�]��{@FG��z9�FAZ��ㅻ�yYA��VX�¢�: ke���T-T�1P��[�@��i>1�g� ��]1��,�#T�4���!��.*��J���q���v���j2c��ZBU��K�:�{�E����ҝP[P�Q;��`l��͛�	>��Ĉ!v�
1N(�X���1��
��j���_�S/~h�E�|�@�v�/)Ea�{@]E��܆��!�R��G����M��>�޴,�����;g�f���V୤aSK��u��ɛ���<k�h�b��2� �eo;���Pfsө���2�]-��$ �B������j��p;5�H"|��Up�&3��ђ^�����ܴ��Ƨ!n��03�b4>N���� �!D�UܝD�'o�:�J5�;�t�A���Ý��[3�a߅���'i������d�U7�.g�WIEg9p�5��V0����3B�gY8�X���}� !��8*mP�Y��ȨP,?��	�1���Z� �gcT�<<�Rw�Y�K$��g.y�������0��)\y��7	(�/7�z�M}��ES'��Ŕ�C�F�@q3(��}�M"��OLG���_��E�h�
��D��Z�ҽ��I�gN]�LlHI�
��<oĠ��'�FNҏ�$06�T�s�Bݤ2r�[剔xJ��$��6B�:i;�mg��k%H���w�t�'����ěuov=G�?;3�'�#�9���r�t�������#�$�?�>��{J��ajֳ����A��3�G���y�,�S�i)!,V�7�JQ-2�}��X�y��P5<A��#T�A��χ� ��Us�8I��=i��Ju�c�}:o� o��ZEܛ_}�`�	#�=[�����+-s��:��,�>�P��)��!���Y���|2��~K8�ҳő:�w�4���;
��5&�e	{z�;{n:&���ZV�Т��K������k�#�`�Z��GTb��lU�m2@/�g��m�cY^@$�%`2�d������Ir�`j�E :� �\@�h�Q�bz�H�/�m��US��%�����B��5��Ma54���&cjjB#�ïfۓ�%��2�[��7,Vdľ`c�s�W1�|3�$>#�.	�E��V7�� �u� ?+11Η��l���=����Z��y�8�t��c�^��ư�k�����8N��F�·���#ˍ���s!1��!�|�b������ w�Y.�N�jI���B_L[�Q.b�
���P ����Q�	�IK��d
���,�qC.ɫ}_Ui���hיNND�7��f�	ʧ�����ӕ�7O���t�S�NN���? 1��!����G ǃ�Zn͎��If�돟�����:�	�5��'"a��zk�>�$��1C���a�@ ��ژ�q7k��i'����ϘG��r�IZ�WJ��ۯ�Gg~狀����E��Y���3��3���"�0�mj ��4ӟXI�(��Q9d�U��K�`��çqc�NG�F�&@��S\�8�Xb�%�l�9��Vg=n�>s�O	$m^]ЩYМ�҅���O�����<?�G���Fڢ%|�Gv���!�OC#�-���FË_+�������٩?��!%.���~&�}����6���Ug���6P=�F����%����/z�<b�a!���K�%��"��\�C5�����q��o�j]\����v"C�I��[M���唓�P�sʻ��d+� ���K�ܰ{�#u!�m'I�R;�{�i\~�< 0Q�� R6ǽ�v���u�F���!�y5���_dj�۾}�!ꙙOPje�(���}O:��i��:�;l�yt9>��D���ƒ����t�o�A�����p��y��w���hx+`��P����]��9R�GC�JS�q醼���!�<�J����?�T�[�x�=����C/$��_\�EU�t�1�oF�$j����������p �Y�&�OC�Jd4cq��ql�����ŅEL�G�t���y���>kX.���A�N ��7*��u0ɥ3�k�.aq��	��Z���hKe�Sv�� ��*�e�����B^l��<N�&d�V�X�W�����n촤1�0��j�/2ɝQ5ÀD�l�?l��ۇu� ��T�QU�	��Ȯ�, �B�*��T��_\��q���<�X��i�)Y3yǴ�E�.�T�fn`�Ou��SB/��,����g5lRI�����a��XB���e�AZ��:�j��L9��a2B�п��=6O5Z�!o68�����B3��rZ��NY���0���[K���Dq����w��"���cg�!��gϽ@�Ȯ�5�B[A��'v�=oq��0[}͟J^����2�!� N�1(��<P�O`�%��9�i�V�`�\j�4��@�_=�߳i��9"������'�
��چ�=�O�ޗv!��PԠ���oi����v�1�q?�r����k(8����&M��*W�A���o�
����m|w/�b :p*�Sͪ,��^m� x��u+;�Ͱ^7�q�[�é���#�?Cڣ-�C)�ßC����c>.��S6?O�?-sKL
�ܛ��u�#���6 �.^�חşi|�5��r���&g��O�hOr�6Է]��}+�P��,}=���L
��wƦ����+{}u�ʖ~
���o��Қl�a�LGq���m0 N��K6�,�b��ȲZ;�� �V�̏��hsn�`5��Y�JU��۬����)�J����3�^X|*�b�����x��3�����<Ur�P8�N�Y7�İ�R	�A���9F�\�]���eן�bo�t��N��p�oRA�l�%�(�f��DR]�G �|�L5�~Otu�@���k�)X��v�
��?��;�+�
ڽC�B�抚3����<&|��UT5]�]�ȉ��:<�<���?��*�<�mS9��gh�5���q�3Kdq6F�1��i��&��Z�#��i���r��H��*��N���1�М���)�0�U�f��vKi�B���x\�6���h[V��Ƴ�}%0#��q�M�1�&�&�ݜ��Q�����քv��'WsY��Ͻ�cʶ� ��җ�̏X�i�+x�W�;'t�ٚI�n��>1��s7��-�Z��I�_hA��[����]#�sY__��=Ѝ�2��Al̔6:�_/�#9EC~Q��34f�wg�']W�Q(����v������*,�/O�46E Ob�\�I9�Ǥ�o�0D�{�ϡ]ХP���^v!�/hu��w]�?@�"���U��Z:�k���YHQF����!h/h,�{�4Zk �b�����$Ȼ��c��Sd3��!�- �ass����ʵ�֞�9��VpJ�WY�ص�T�BL�{�b�5��<:o���	'��N��D�,EZ�z4p�^�d�m|���Q�z_,\+���:�1gH�/��O�wMτ�Em����ֱu��@e'���iYέ"Q����Ki�K?���x�>���C�ܴ0G�`1���|���>L4vz�;s���aw��^����_��8p�\�~xc�[�(OТ!թ���?��-�סgT4�^O����ή���O�_���X*O�V��%^ur+?/�l��˼P��g?'ضͩ�@L�o���D6�=x�K?y�1��T%���x�@��9LU��������b�������T�I����,y��[{D�Ճ��f${Տ�U�QNgi�#�'^�r�bK��x{_�H����u�:t��(����,�x]��x��J�h��b�
;V�}I�H�H�1��G����*���m�Hq��/TS����(��'��6ݟ3R#��O��!//�E�����iKx�Գ9�P�i���.�.'����x|Qz�F���v��Ǔ�V�V)�}y�/HJ�u�I-5���A���dNp��CRܓw
E��-Ѓ���bx*�<���~�g�U={���cd ��j��߅h��O��I�_���#� ��2�`S#[�0��� �Qt�`�l� ���P�6r����R��
�0�wѽ�L�j��n~d�x�,��ݻ*[<�&F]�oth6�E�}�q@�jMC��f���<��[�N��=֝?��s�"b�h=�i�e}��z��ǫI.6j��6��%��k�)4��yԄ�<[m�?�1�$��h^��qK��}�����S�ED�-bo��ƥx�����QT���ǳ����JW�X���˭�,~C�� H#M��:ςĸQ�``n��꿿 o��e�lK{S���J���x�#�#UϦ�Օ�� ���cc��/�S��Ĵ�~y����t昼�@�l:MfC�s�#�0QР��K�I����G��q���#"?$�������Aﴌo���ԇ;��Ƌ��Ѐk�ؿ�;*4�z�e����ŧ*(�,x��`�S'�[2}���W�Q�@S#F"OTK ��i��P�f0?��E�,;�oާn*>�@�ٗ�Sg�)�����-�%�^	�9ȚFc!|���+���V���3]���q� �m�9~��)y�d	'vvAc�{�ha�Jo�`{��2�\�N�ڪ}�,�ڳ �v�q��r!�B].�u%gK��P�����%^�ۤ����0��I�j�*��K����5�*���L�*��+�o_����T�!��?�:��W7��6�S�&��r��|(`�6-���u_��:8R��8*n�5�v��V�"q�'솬]D�����܅�f���!滙�?]�������� L��V�/��'3t��3�I�R�"�JCI�g�?�:�m|��X#H����0���(p@�`.�pµ�B썙�T�0U��������/{�j�7j�8l�T �@�r��.'oC�,�
ᣒeD��o�3�b6��,e���w���
`	��+��êx� y�E߯�xm����ʅ�>~I�W��?P�MAf�@�aE��
��v�k�uO	Ӭ�Z‗���vɖ	����ݓ���z3�um��4)�|E�T��C���r�&�� R'(��c�Wz4���!E�D����J7a����S����c ��OK�Vv�~Xe���'�*k8�4�q��bF���R������Ԭ
�����trGgS���mk�y�߻��^�&#�����d��D~x�H����CdX��-4�N�(Q�~�R�H�E�)?��{t�T�Ƀ	Z�(�e��49�)&SH��ak�UHc�9�u�e����3$6�3���GD`e��b�V�v�qЦdߋu�ԍ�WS^��8Bv��x�[���UE��?�Rk����_�k�(���F�4�����P=z&9���D�n��4$h���}B��'�E����K�
��)�14��]IO}0�,�	x��Lnt���a�r�V(�D��7�*D���1,ĒN�7�O��R���[�>w��a��W/HY��/$K����0"�s��jw� �r�)G���fu��mD%����I�&��Y]RvQ�ttۏ��n�7A��(�`sY�B�X!��O���s�ɴD�b�І	���}�*�G���
[�$����堅aZt��k
[ħ+��|�F_B\�?��P�ݹPե�l�<�S�m�6��|�����H�F��:�f"=q�{�B;���1�x$����EL6h+f|^�	 �~@^��Mn���NftQ"���/�%�%g�,�[}5�Z��3�Q�Zj���W��[l�L�7�q�"���\ĶѰ{&����+[}a+����t�*P�<������W��M7�ge3QT��G�%k����Ɏ(r�T��s�Uɳ�<� (�����[%�zu�-q��X�h��n�k��[tk�?"h�ތ�-=�x���)���,��V��Xz�T����
�g�{�=�v��gh�-�{���'ư׉���a�&_FD��Fc��|���}L�Nn>�g)<˷_�=�LIq\�~������K�E��`>^���gȻ�m���M=�2>�>��(h��*���QTx�僛_
m%��_����M���I^qR[��b=�0+����}k^�j\Q2@+Lk9�}�@*'��35�'J�9�V������k�8	�����Uc6p�PdC���!b�ȅ�z/��A���8A��=����@B?v(�I�X{��t�����&�[v?����JLp(9��ӷ�ۗ�D��6�7j;���)�_VC��of��Y���c�߸`����8!��b�4ۛ ��3�,*���!�l钔����z�����r���i��{�3�P�睺Ꮘ�qZ��c�[8ZC��j�&�����a��D$Ư��~7�Q=G��ٻ��n�/��e��z���0�Ep]I�T?m�}�)��.��ɳ�Y�s@�*�qYq>�L�~+�������3Q�ʓ=��a�������b#�W����9&ƍ%����>���'��.+\� 5��/�{���[��'8�Mowh�1���+�	�=Y����j�1�2�w,ʰ����������E4v7Ht	$�U����!<d�=c�,��@�v���'�;{�c:��y4{q�,���OjV�*HA��_@0d�����~dAs�F�F�M՘·����|����׆��z7Lv�ۃc�	�З���ݟ����!~C�J�2�)�j�d0������Na�n��r�^��x��
| ^��nΕ�?s���#-W��=7M�2E��W1��ڍgB��F� �HjG���.���qOzLp"qя%�B��v����x����l+�G�4�qe�ڎ��������ˇڎ
�9����0X�IQ;S��ۛF��to7ohe��fL�5�[���D�c�����ø����Ң�Ȑ*�c���;�UM�;U<�x�maG.Sj��8Y�ԇjؒ�t�/��W�b9e�1=���z5#��,-˜,��1������$���NR��5�����W��)�ٽ��ꁖ��v� ��;��Ѣy��E=6�+����&xb�9fmw��`7�}�󺨮½e��V
0�WrE"�����!w-�ϊz�LN�F�>�#�|��є3a*� e��J53\�ZJG��W�JQ��9��n�Pcm
%��>�X=]����> ��b��vz@����!�V�E�}�8��UЙ;
-��`X�ѕ5tW�z^ï�TU!"~$'ߡ�\�Y���Z��3�3�|��A�>�ߪz���L�I��
� �L��� �|��,����(v8��V<����K�Aȱ��h�.x0���ڒw���5G��)���|`��i�e�*`)��ȅ��fe�f��W4IG����6��o�c���%P�P���r^D"s��#�@��[Q�.HA.��eh��������L�g@u��vQ7������s�oo=P�)�86L��0\��|A2UK.�����5]���vL5��(�r��"|;��S�% ��<���_�����D=߳b�Do�W��+�Aa,}I�cwam���mա��;^�&�� �@&����S���Y�^��:칋]r�t�݇5?#�L�|���
�4�,C2X��"�f��.���ܕ'�Gv7%��c^Q�L]�@�FWc&c�m�5�����3���8b[l��'
b#���׷�ZI���1�E�_iZܫ�,�A�g�SVNӮ:Ux�B��,ˤ	��T�f�vHEP�(:䐟to���Q.�.g_�W,Dρͱ��чWę=��P�9��2)�~;�0��֖�8ت�� ^�+4��s����x���K�X��%�!ED�Ɲ������-2�mHHl�����Sδ��{p�E�����_Ж�����IEh:��'��i�C~{��//���3��a'��_�m�6'��x���k�I�J|��,	Tā��b��R�E�S~w)P�Am�'���>���q� ϶k�٩�Ka�J��V�O��0���t�G(�r�0� ����H�
:�n?EMF�2�n�ӽ�r�������|�~9�fR�~�uf�#��ȣ��KYq�-�^�c*b�����^�Z۠�t��P�W���U��ך�s��c��>EU���_��.Fb�������l��s8�R%�ly2'��$���F.� ��p���S��p+�e��o��@ �|)|l F�Sfr��>u~A���/,s�W��*�a��T*0��{�U�����r�;9\#��~&�s�[���;���u������8
]U���ر�}w���E-&,J�2�����ڷj�@�`i�d�ӖHaq�T��[��*.U.U��LQdM�
^+�g�c�U�6w�q,D��+D)E8+59��P��