��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ���\::��_5x'��n����%A*/�Kt���D6�O#d�h���y���6g�����=|g�p��X.ftk.������ُf���0 ��u�A�$.?c�En}��%�9�H"S��������Sg)'d��B�f��ꎗ��"��,ټНea鏨�꯷H�f=���^�/�p�Z��RAT����:T�2s��q1�-M��C����9Ẅ�(��H��Z7�G9�d�����v�]Ȇ{��?����Es�{I5�f�#\.�=P���.>���T����Z����t��6o����ܦ .�3-#�I�k?Q��#�h;�E�
ڜr�)-�!_V��y).U�D��qZ�0���Y�BA;X{x1���Ռ[O{
$(�[�C=������XK]V�,�wj8���V���ee�S�a����e�rBV!��;��?�ee����T��S����N����rf>%n�<�i᫈�~�Z�Ǻ�xT;�ۜסf!����a7.*���g�����@�U��(A{�B����~鸟��A�I�[�yV�U��2��v�J��O*�6��eD��^�F�L�N�=���#9v׻�Lv��V�ϣa�� )��
h���j\�\�ڀ�G@k�"�=݁�%K��T"�*|[��I�(Iئ�E�o��ۗO��d���8�mk��.���V�H����uP8)���8��V����6�:�ڰ�9$�"�
~@_��fs�B|���K�+���澥q�f�L"t2�_��Q�-m���N���x*��`��A?G!��zvQ vJ�h]��.�$��_�{d����(��a�ԛ�tGM��[5��P�RG���J�0��I�X��ǽT9��P�� �Yl�����JS��,Q2�j�r�`UWK�E��ϳ��,VZ� �ko5}�I�d�tg���h_:��Q�����L�w�7�Z�DQװw���C��7�S-����\���f�.y.�V¡՜��TU0b��V�V�^�}iO��je�+�Ih�C Ȣ���m����3D����b��5�z%W�À� ��ЃpZ#
s��ն�`�"�D�{Ǻ� �*��g��8C�_�!^S�m���˻_5����wz!�OH�دME�����c"��!\`|��9�g�k�[��%Fqh�#(��7_r@%�0nT���SB뛜�I@1�kd�톿_x,
/5�~Ñ9'��f��"����{�����ϗ����%/����	�3 4����^�T�O��%TXj`�!6*GQ�K�Ab\CyO���R��䍶K���:$��?x� I��8?:�G8����mƱ�e��x�CN��ĉ�d'6~Q����P8�C�1IF<�$�{e{]����.���Hc�"��!?��R��t��r-���'�-5�~hF�ư8�e&�n�ɿ菒Tx#�j���
���e�L�
�v�Dx�dMƥO;�F���o��؏$*��[��j�+�����N����[ˡ�z� ˈy75�i������W�$���N���xf@lЙ]�����G!�0˸e���G��g|�J[������2��z�8P_1�L��?m"�L%仔%�/`�N�s�����(�q�U��x�d�V���f� ޵
����}�n��0�&EL�	0�R���5�y���n$�`�k2��\l�ӂ��Dke-S�ɲ��$e����~��r���ѻn�����i�!ش5�GF�o� �&V�!i��\���5ͳkب^fH����Z�`�u0����57j5C������ts3��g吳)�� ��m iN�-�:��C����ʻh5M����g$�:ɷ-�T�Vf�I��+�pNgρ�UN�o�PS�w� y��g���� �b@  �5k ��:d8"����	�J�F���@n9PiS��H��$+�$%'>{[eT?���af���i������:z�o��d�,���>����I�ѰF'^K�S���N{�櫖�A��.M5���R0
|���jx�����I��ޥy���L��{�U�����3����sD��s����~�n�u;#��� O�1`"U0�^�z��(|�9^�Qv�\6�X��h�(~�Ҝ3��^P�NV�ދ5"����1B�( ��P<�5�ʤh�!���n7>GUαJ�9>�M���x���	��.�P�"r�!��X��1h��~UnHb�p�lm�tTX�G�eO�����-��k#&or̳�ql�N���P��_9��q�>��r���1�f1�4�C��^��UW��L����fQu�����~#>M_�V��f�/����[��F.�|�b:U�Ô���|q��o���0ޒF�I�	� =K��oJY��B����Kze$��Ecu}U��oq����L9N3D���S�,��n6K��Gg��>�*W[;�t&t�Yz�Bu��+����~��-	W��;g����y~�F1��6ypM�d�VR~�V7�N���r�[��a*��W���5����<q#
"�Τ���(�����B.�񫔰	s��8��G-W5�?v�,���2N����S����e�T����7��8�Q��Z4�Y�m����ڌ�{�߀Q;��Fo�J���s�q����5�]Me�T)�``���o�K֑F۰�NG���� E������V2�H	���b�5�0���p�7ɍH
ܰ�%g��|U�U���P8���t�9�/��C2�c�kGDE�0������8�+����D������+�&t��3U>��tO*��L�~���%�+2�=Ka�A�K�'~�O>=�����	�<��$�å��l�6&��Vp�����?� �*t�W��({M��"�M��-d��#� 08ë�.�����C��BFEs�`1�G���2f�����e���)�\�X��5��U)]T�� ���.�(�2��4�U�ގ����.`%r�����^v_�0��l_�?��0?Z_l^�Q<�}��^�A�ňϏ�=k�vZͧ��bʱ}=9^	���k`�'J �.q�T
�T�e�i4S��M���['�V&ld��Hy>�J[����u���#��w�
u��cB� �;���A�D�&�@8'��V�lw��fK��D�|��q�0�2*+i����7�g/��I��B@��늱/ns��?�P*��)�h�>G�xb��ߜ|G�
J��0���V�7{��Ö.t�E?l� �`'�88���ƶ�<f���竺�N�=e��U�b%w���j�[6�d����An��]Ll`���<� �	T�k��m��|y���xɌb�\]�F%}�bd��h��/�4'�pn"���J
�$���j�3o�P^�W̡S���t{���D�1e������G�5}Sb3���:�~L�
n�F �?{ģU�L�ol�:��Y�	���:���9ӿ�J�?�^eu��q���զ�AZ �xl$�>�S�&S��ǯ�W���1FB�Dɫ��l%�"��8�a�;�YɁ{Q��ʨ&3���6���<Ld%y�uژ�;[�}��z��i7>�U����)!E�ˡ[��}���(+<i�y-q��Г�����ɚ��m��$h��b�|߆�;�ڦ$K�]�i{[6���|8x��_����
��|i4P�r�BCW�?ؓf|R.�O{�YZ]3u�z}����h��v ��7�;���s<�X߿���j�آޣ�l��t�'�(?�ȇ^��@��ax���/_��̵�̔i�(������4Jy�3`@����mo�ν"����ݩ���V3P�)�z����(tif��3F����e���W���uh���W�(���tu�3�NY�ӎ����="}<j�����y�V�y�Jr��j�m�ƌ���
�P�U�q�~|�!e(k=Ga=	|�֦SۣU5��/��<��{ l�4
�u2M�]�6���+�|��E��b[�v����_}f�BGƏ/ �:�L»��XTcq�%��|��1�'R�U��p��΢|����}��������,�/���YU�n��G�q瑖��H����^� ��c����_'g�����t�Wlo����6L/]i��b��U�HV��Nu�t��6N��C#�k�v����^A��w��e�[�H	pX���
���!��۳���Ia�#�T�����ҰXZ��N]C���埊*1T��幔[X_믗cU��& ]Ӣ�~�X�L����Qu1��n<d�z��y�+s�����l/��D��_�	�g��e#�EҼz���n�d�8^��Qe2���{��`�%w (�Xo�x%8L�[���OR���q1��F�O<$a�qZ U�}��Q��ʁY���\�͌�3������_Pj)5%e�d~i��·������'���&Y:,���ձ�b!���G�t��V�����,���Ru#~���h�����"���T�0j˝��a�k����V���۶r��	��"�U���I�=��/%t���̀��P�m��w\����4���3*N�Zt�yE}EVL?Բ�UP)�L��*�=��J�h��i+��m���g���l0V���D��2'!������W��Z!�E�^���
������|ȵ�Ux@�ײmV���@t�CT�y�?�ՙ��m�eqn��pHN��E��×�%�@�+ɶ�q� f	��5d�:5R���od�������yB�����~��F�K��{J�X��5xY�5!|�. �O(ۮQ��ka�7)���j���z��[�SU�C�I��)��� �1K����1
��i�i�����T.x�:����"���CFQ�ֶ)� �~��Vw�Ӽ�oVŗz�����=Y��6�*�ҕ�'��HR�n��m-�ݺ��?UR��K{�!�X�SP�V"��Ͷ�qL�����#��mp��bTa��/9uY��5J_:�ޅ9�w��^y�V.y,ʶ6lw^�[�t�!ܘ��f*���ӣܖ��G�;MJ&�n����rz�T
p���@�[�Ҵ�u&'��8<���td��;n���{����t1����9�
�84��礊Z�=.�(���6n�{N�LZ[��}l�k���r��}�T�I C=�H''�9�-ܖ����AX�nw�.��>�+y�M�r2�<����[m��;m3/W�ҫ����r'tz)J�vIi��c�I<�4J���V<�ڸ(��jV��в0���=`����#�"��>��T{�n�5�����A�@P���X�ڷ.=h���Gt����X��s�����g&�!�'4ɑ�o�v���<eR$�:���{W>ͳxM�\��/���E`��$"ӺIc ��.�CZm<n�v�ͩ��4b$eo
4ӓ��~�4�ꬿ&}8��j;O
�2.6��F	=�S�/N��'l8��:_v�>,�)!�3lRF����"}�!]YPv�师
{�����sޤDp�> Hpdy�x�=������=�+��Vw��0�<�0�&�����g�m��sz��("���85��C��W��$�{�����a"&����MM���0;��K.4�6��.�D6����@D4c��t�&�6���>�?�)����vUp�����'��r�A�K�<����W���4Jc��^/>�&.̕`�8R���v\�	tT�`D5�=%�ʚw�#�n�ގ��K��Ȑ���w��DkQ�?����Ȣ �v��C#q]�+��,Sµ�|9��k��Q�:i%"1�$�a<>M$giJ!'\R����6�ސ`��$޺���L��ma>�&n�|&�ʈN�NB�E5t�tkUk��<mP��C������o�����]&F��Y�У:�)���W=��khR!��-�4|���ó\5�A@���4��?�5�0L:�ю�`�ڡ0��@H,F���񚚾}�(�pi���Ȭ:\��a+�Գ�U�q�,lnv��p��GN	�w��>��u�KG�2+�a��UW�|����Q�хHS=Zɑ�X?�Q�`I;lN��#�� �i�y�Q���^wx��05>�Q$�~n�˱�	A�H��s�`bax����o���S�㜒Π�X�I���$Q��\������#�_3�^��j���Q� �~��JF�i~��� �-��'
������Ha��Z}�2����j��Î�xC�5�1i||��=���b[
"����Z=�Ha�G� �&��}�<1{L���L�(R�%׊0�ނq���W�x��+f��u.�0I�����ތD��A���$$W� �Y�Z?�q
P��e $�������y�
&�r��gF�2v��Hq��%� | 8z�{SY7ɚ���tb���0C��G<��b?�9��F��c��e�w�M�;P���ArA�?#�G�����Ɛ6S���C..NF{�Ba�l�Z�l�m�T�F�����X�|*�{ϋ��U��r3f�Cڿ�Iل0w�7�X"#^��ͺleb5�%��w
 �㪊��8���W��E qV���I���:���@����,OB�?Kk�oΚ<swڮ?����(��� ��+z��9���������h�ؤ���Ծ&m��F�}�T���w��Da�1�}a�PfT���%Rڝ�ox�-�u��h�;���B��%�ך���V���W匜��ܚu\
8�9�E�E�`�]^cf�.b@�A ��b ����^����`�=6w��%�-��l%sd� o�ۂ:�TÐ�A�k��Sp#f�k�$E]�ʡTɇΞG���0Z�!B;�$w�q(�iuXUG"�}ZT%�Td���c!����$�όꂵ;M֫&��ITg;+‭{Y��j��N�`�ѫ���ϘNP���@+��%5
)q�#�+oy/ﵰ�Q��~�s�(�]ʇ�F�S+YWB<�����K��LZy��ƛ��~8�~7/��ZLl����R^���򠰛�KSO�Е� h4�I"���	^�\�����0?�����o�b��y�]�a���~��61�3b�Ǯ$UN�l��!��}��T!�MsU��!~Rɺ��FX'�Z9	���r:P��� ��6 ��FҒk=<�*����<Eu��fCsE�'�"P����0w������I{>Q2�Ҡ�n�����:.a�-6����￱��.2N���I�΀CU�y��W+��Ɓ<�u������Z�^)�	}~U�h���hWc��D#k@>�z�I�9@O�q���M|RT) "y����{Y��Q �E�?���1�7���λ���8����DS�Gi^�����-���1V'�U�%�8&�ο��r����n�nd^m���C>W{[���С�����o�����m�W�=(��ڒ��)zΤ� �+� vu����7��D�h|jh��G�̦9���1j)��ԡ�q%�Rlp�hOl~i�U�@$�bM2�u,��=�ʲe)uC<�|������0� �ii� �~C�{�l,YB��`�$�4p�ğ�Xt��u�I�u����s�.� ��~\���oW�dQe���["��vM�X��Mw�nUFW�'�f�5�����M�W(��q��ڎ�y�T��i�:�*�1*ڻ��vPK�nS���La�E�Aʇ���%�n�*_U��_��"<ɕv��
O�+(�fC�/�e�c.o[��V�6�����|��΍���XO�t�A��o]��*4�k<�z�6T�N?������\�3����:z-ھ8���@���]=BK�_a��?����Y^�-r��䆄���G���fl�Ԗi�]P�&,H~�M����q:�!=v(�X��C� �ڔ�ҟ��r����֥�_�X�e����F�V)Kr�-�X���%[����V�������h�hVXd7�P$�K���px�/ܴ�9F�&�	��(=��Y��p���퓾؛;����������(�:���fx�`�Ĕ�?k�/��5�����9MS�6���Vx��u]rL��})��IY��DU\�"Y%�mP�z8-��}@a����KYE�a�у��J��2<��l���C܌��\�y�w��r�{�ĩ$H{K�����Ʃq_we�����;��Nb��~����	d���d���ۀ�B7a���^J	�L/�v`��{��)Vs>�ͺ!az_�_�W�H�a�"d�W�o$ԖL�Y�� A4ߪ��SCh�Q�5��e���V�Ԗi@��T$i�]y�3�V�w�ol w���μx!�Pu��;S�ۣ�53�1(�W�9��	?�Lͩ�G6)��WJ�PS��L=ֵ���0��]�z2�3�Y}ʭgш���o|v+[�qu�N,5�n�l�d��H�_��:��p�ʃ��|�����~o��B����?4`k�X4�}kG����B�[T�s������H�L�-��B�)G�������1n���N�>Q9����o�����Ƣ��\A��}�e'�t5#��!\:����sz��^ċg!�6�Y�P�v�p6 �uMdz!��C��+�y�)6R����t��	/M\���E$nB�i��#m�}�GPD����s!L��דsq��`�=R�o��V��"��M�(Z� �鵌�+������t؊0cE��q̞ Yɗ����!c<D�x�Eܸ�4&�ШcpVy\m`���o�##��wUc�׹i�$�m?�S�GJe���=�}�hs�(���ZH,_��������N��\GWбө����V3��	�d����ٷ
�Mf�,=^��J�ࠅu�k�q�<*��_�MW5��0aRb�����em�~��%�B�R�e���'�w�U+���pJ��H��tj@��,�,�Ӻ��j�:�-�,q�C�<��k�w􂏅���qA%�%��������ވ�Y�V�m��S�6sd�����Z�t�@�B_w�f�������;�� �e���F)i6n�~���(a�>F�*�,��.fV]�x��=��1ap��	s���Rae���ӋZ��0@_�)�E���p^��7�s`1IM�\7��)O�}��xQ�:� ��K},�g%R�҄|�u�����f	Y�e^�v<��$���EÖ�P��z�uB1s���'�)L�/-���j�4�>a��2
��o��H]���ݸ]��y���z�!����������&����߷=K1�]@���r�߸���ڭ���`t�%�W�G�[�]!��x�$S���3��k"�k�m���u�Y�4�R*m���1�'��˺���R�����4�
���F�*O9P����y�7����#�� ����7����s�t��4����-u�,�-[vR�����w��a��8j�!�3/�2�,�X���b�+k@���8�r3�k� �Ķ����Cd��5^�J���._q��/f�z@#M�I�b,*�u��u���c$@���"��N�!��p��g��t��Hi�Z��X-��sU8�X\,�P�q��bA!T�Gر֕A���[n�3�c�d�N��KՏmmz-���d�Ԛc��#�
c�5�&E���ޥz�E�~oއ0���0!���E�p۪�����w�m��z��1mR�l0^��� ��3t��2g�|�����v,ŷ�0�
!1�@N�(���{�؍m���J]�vj�@z�K\�18cV3�K�y��/g��f�E�|�{ݗH]��ʰ`<�g�c��-9i��Q/c)�N�g-�����G��rp�W���lI�1�^߯֟~y�ػf���ȉ��3-� Z��H��1Zp63���i�����T�������A�j��d��B���c��~4�������P}��K�zlZDu��h�˙Fl��בN�M���\5�[� g�@��?X�n�k�����(o���H������(-����j'5�V��R���됑������ͤ C.��q� G:�K�V�A
��j��(AI@F�ųCF"�ߗ�(�B���W����(�q�ó�8���2�g7�71��Q b���U	��g0si��wgt>��]�d��n>�#���ۼY�r�T�������_���gH���?2����l�V��{����t)���֕��r�d(�����ި��̅��y8�n|b"	U��髣q�� ���֩�P��X]��r�$m��;�}0Ԇ�Z2!�.��/���2e=��� /+!>$�#H�d��,~�jL�P*���G�O��Cd�+5���C�<T�8(�g�#,g:��-�0�������{�[���<ō�=��Ѵkf�4r����p<��j�(:�f��(B�j����n���+���C�d�!F��R������4ɼ��1�7"' P��Eە��G���HZ,<��b���>�  @��t7BY����t�˛�`��ձ�[aڬ#����ԙ��$�E��c <����깏�3�?`�La��|��N�U~`ء�r�-Y��F�I���ݸ���!��N;o��}�<�<�,6�=cL��ݢg(9�r�g��rC�?ن��l����� C���^I����6\X������歨�٢Ә)��p+�ڋB(�7�4��\1F� �7=�Ix���Y�bI�O/����rV�_x��Lz����,�C<s3�	IA��Y����i��^����],wb�,�=j�Eؖ"Q�n��{�祾Ζvb�E���R���Obo�(Ƈ�n�U�`
ou�<w�����/�i���ϗ��j����K?D���Q(�u �fu0w��!�=h�r�e���(W���L�O��+�M�z���G*9<����)�"?�[�=8��P}�jL�5�a�ٙ)ȃ�i��u^K*c�~�2�?�	�h S#���'z�������]�Gacg.a��@�+X�C	0�������!�2Z�Y��a�bՍ�%��U�IÀ�)TۏA%y^Lq����4�_�ť-] ���_�ϻ���n�R-~?���h(���^��W��0���m+���?~]7���U�5ݿ2���3MƤ������t?�sjr��j���ń/�B�d�9L�8��{F��
�
E��	ZqN��X��(`��D�}�ms�L�`)�}�A����-�޻}�w*׀� �]o_&�$c���W����(fx�h��&�ʾ@��n�u�Ur�<=���Q!�u)�����y����[h�ףp���6��Nqa\�kI��pEUbZ�2�0	�7�Ҕ!�RY�Ǽ���z��,�*A�ԏ]�����w�$:^|�vyDOw��;�/2PX�z&�7��pot��=�	��eX����D�lE#����=G!��)����M�i^0dr`��L�h�֣%nU����tz42�����[>f6�~T���UI��hm��m��_�C�<_ɩMO���Q6�H,{��H�����UQGA�=�3�=N�����^��.ͧ��_�mXU��XH�ؠ�hA.�%���&�Oߦ36R���p�7%��野�7۴w�%�I�����Ɋi�
񝒶�J�zH�©�߫�L@\����������%�qS.���H�W�g��ǚ���M�,�%�ߋ�eMl�P���9M2\SOz�B���/; Y='�Z��K��\4_�' �S̔���R��9�Ky������c�N��zc�M���-g�X@=�$]���N�;�=S5��an��@UȮt�^NsX%u4Yu)���T�Y]�`�ǌzx�N����'�SV�s�S	�VИ��x�1����u�ɩ�_8��|����Ρ�[�.2�����8��o���Q-���%�+r��l������1�Q  ]�=��C�s�8Fr�T]J���i���n>�,�M���\�J���O�����u�(���ݲ��p�(\�b��[�W��`pͅ]����6/��T4:���#z�ؒ{u;D�	�C��:��97�(EY�.l���f����֏8��-J��@P>g�(u�S�n�Ī�s��c��5w������đ�L;i��@��`E
���U�[Y��E�����xe�7�W��;��}� |Hϡw�y:$
�f�S���@%���wG�&����K���Sͻ��kݰL|ՖdZ��������UFuh@����+`��~tF��"��Z��q�h*����J��yU����xm�}����팶f��[1H�'Z��+o�B?�q�%�sa��:��H*Anl�`ckg��=��'A�Ʉ��c�b��mPwGҬ�ڌNI����{�e��R&XԱ4R} 5�Ց2�:ħ�4�w��V+Z�����aK���E��B8O�����:� ag~�PjV��������F�]	�yԐA�u���OʙPA�Q�v͕��-�� )v�ur�;��&�*���
�g�W��V�n��ÊE����;)�	Y�E�O��ZQ�����)~
=b�4�&h�N/�%��X<d)��(���ݍ�F[zT΁9���0J�o%m���8��䙳�� �U�cZ/��@V7��hA�H���`ԋ�.a�hR�:��Ú������J��+�{��yq��뫟o���>�;��$-o^{�<h����:ی{o"2��!<?R�Zv��xf���� Kf�f�^���¾B�ȣ��=��ZuՒ	��e����T�~���tlb�Z���fI�c'|]��$qۏg>_������`�~��l�Ț���J?+&	�٦�T�rES��=���t�g�*i�N+ے©�n�����pY��:Zk�F�܀�h��@����_�Z����+���J䬿�f�*�B�����V�G��e��������F�4E<����m�L��a�5�� BK'N�S�������g��1��Ը}��n,ϕ
� BoW�0�U&��*�����*�f%��Qm��/��+SP.���w�/og�c���.�=�_\�L�y��Ƭ��[�� �"��v�)�?>��Q���3O��%��~h�n����E6�����1=+�G�w�zU�uc��;�ZY��sJ��¯���QΧ魖�D�
vn��f[��5q�؃h+7=�0dXĆ.u��Z���<�˳&zBr�f��x���G����$��45[��	�o�rE�N⊚�	z`5�J�d>,+�B��	l�+$0�������WX���2��fȕą���[Q�Ai|)�hÊ����R�&��S��st礴�·{�� �i��4�ȧn=s�g�>O�v�aw��������A�����e��I_�y(�y�}v��	��>i<-��A�I�?��R;T�������qK�{f�3�a6��p�k^?ܡ����M�VT\������SKY��_�x��o�m�q;��?o�C�ȱ&��0���P����G2S����{���١��HiW�rm���H��{���J��'��y�1]�!���Y�H��V� �c�;��(�\������Yw�vc)E���{�|���;X�17���\�� H%Xb��W�{�M�P ����*���J�+9�I�4�ǫ-��qW�/�?3�����Fl��0�w�\���1o����Ԇ�E�dM���[!5�nH�,'Äh��ߒ7�3c	Nm���	�l3&���X������8!-���}I�G��:�����gi�3��O,ˑ*�^���Ŕ-Ȭ����ߢlzyS�d��$?$)bx\2��C<ԛ'!P눐f�{6%�J�t �s`.o	���{ҳ)f(��@+Ҟ�1����K��W{P-fD�0Ϲ��`=ta  ������r��j�����ZdV�^�=\�� 1?u���.{T@h)��Y�<����9\�Us��j(辏��^�ȆT�:���r���zO�a1��.�y *��v�lWm�T��2�xaa~��p�M�;���P�Y�3��Om����e̐�د])ւ����j��*ykYf6�R�*�����,Îv8�af��ָ|DFD|��X?�6�Hmm�N0ǻ�)uy�
�
[��3���w�:�ތ��mP�>E�;~�ڱ�xK���JΖ�II���ji6T{���� X��\���A�Z2(U�A<aY�K�ibN����O
[b5�9�`��:�E�S���3���،�����ǡ�u����}}��d��Jق���������v�S�}�����
����Q�Hn�@�{AQڙ4��;b}L�@����(��j�c��տ��a��G�53��J�|J�d%?V ��ݨo��؎MB�m��P�
d�+��^pnR�FA��A5�aY��T���@Б����ip����z�a����]O J��(��7��k��R4J��D�d���<l�[�w��$�t�鰯7^S�Cn�J.��R,�s�f�����(X,-��'H�[�,�b�
Kn~��ta�E���G���c�2�b��Nfdn@�GH�d:#�xO�Бg_��3	6Jpl����Yi�h��\�*�E!vd�'$A+h��.��:U����m��|�t����ʹ�s����s���G9��	-1��Μ�a�xo�9�Ps�O��*�iU��A�]��)PX�+��_�<
8P��:\�R��Dmn� U�Dē�跽�n��g�B �/�K�Jj��ٍ4n0������LTz�W\���bq˷�e$XT~y�I����O�<[O�Y�Q.��n���:��ne�@Zo
���&x�F��՞�.Q�S�(�`8��`,�n�A�b���,��W�#y��x����"���!>K��{�#�W�t[W��������w�fH	�
�J�L:T!��)T��9��yn����5�a��r��5�Kw��{�s�̋m��ӟ�s-��d�(z�8-�&���i��&֨��M~��G<��d>a�b��="�cx�EL45/ �9-x���b�z���ѥ�S�2�,��Y|��@⅁��1g����r��&��ӐO����6b������'���J�A��>��E[�gj#[쯑4���T��3Ё��#	�\�-��.��;D��:�A�0�|p���f�>��jn����H�ځ�l��<�d]���I��@�}ɀo��5�|̈%��D�B��?�D�V���Ț\���܋�q4� _�)���k��Б+!���T�TȚb9K��Y�W�D".ȟ�TJ�����,���0V��kI�]荱�0��EVV����R�¹c���2!!�-���f�v=Gp+>=�qAx]������W���M�u�gZCor'�֥~+����!D�b���%���	�^��T�(�us��ul��(�R��>Ǡ�ٚ����q0�xY���&+$E��|�i��N9Hx䪩�3I��X�p�qf��""(ڝ�.����j @��J�%X�G�P�����E����-MkO&����}�d�2��C�B> �~��@��R�+��+���J�z�/�Q�K���0�A��MZ?��3��W�X{t�eZ��v�Z��t6��N���N��1&�cڐ���BvR�p(��r-��Q��i*�5ٗ�$��ԩg��k4�!A�E�|���s��"t��[gRi5T�3x>���|�4�Є� 5��\�V�O��
��#����<)]�JB�3�ol����?A[C4!����DZ{���q�ed����,O~���D�+��t>�R)e_yXz=��	8I����	Ӿ�L��2a�T���03��:1l�gu��_w�*�y$���v&�Q[t#�܀�[�6��ł^�Bf�҂L�F#�S����`5sR	 ����s7��A��	�ݫu�&�ɹ��m���n#nK��j���xq<Ȟ����1Z�,ȹ��m��}^fХ�����W,Ŋ����	B's�XK��6�g��gB&���:�>��%w�e�=ePf�l�+C}c��a�qɦ͜	/3��3}@	o�*�o���ќaCN�$����7:�喂�m�.�b �.��N �����dq�_v�z#�3�{k�n� ��Sco�ݢ��2�}L!C��nr4-ʹKP-d�� �3�m��� ��[6(�g��4�ˁɈ���A{=j�*��ٺ^����%�a�EU����H��"a�ؐ5�A�t������rc�2�E"�;H.~@$*(@^��h��X���Bj='L�/��p�~�׫�-�d��;�]?WTb��΁��}U-�%�tf��P҆���Z���Ro|�?z��s�9<����HlFJu��E��E̥w�F ���0Ɇ�;g�b^,�D(�u��^���	7�{�rmj&�aԝ��V��ԕ�q�2�:�|Z�o������V�!�0��KS���k����=$Z%��d�yP57��|��^�J:$���ŪV|>�M�*/.�4���eP����S�5(л2�s�>�����=@�uR2"թ�'� ��Y�G��U�HOM�������/�m�&4�� ��|���c^������v���G=�X�̬ռ� ���M���v�f�,��) �<��;�M����d���\�{�q��/a�����^�w�&�g	b�v��z`���D^�q��0?� �a��r����j]�!�cR��9�x$7lS���Tk�}{#ٺ�|�g'd:eߚ�@���b������@�#@|�䁫6�m�X�U�2S���	}Sk\�Nԡ�`UԒē;�ɋ$��6�s�{�$gY+!'�ܭb��,��x��p	���'s��~ҋF�O�y<PG����>�iXGo�i�G�g@2��&�2���0#u	<}VB�:��z�Q�����w� -m��R�����2��<��g;^R�lI��%Y�)�e��'�U[�
�#X?O9G�z�Ee�I��(c�K�����GC���f��ǎf*�f.��m[��/��:����Rf+"fsn�}��]u�H�.���=��=tM"��tbl���?�����zÂ�)Q|W�#9��*� ��Lf�k!��6���7K��z䁹U�>I�Ȣ�>���-M
�W}_$Z6=?��[esm��oN\`�vU�����xw�x�S{v��cM}�H@��$ٻ!�զۮ^��w'k�K�1�;�q{Y�1n5������y�����#8�v�8�~�d(�]Ma��
�D7��<�`}�t��}q�-0+~�mH$��mnIð3�0E��Q����O?�r
[���0�>�2v���&�ݢH���x���w���Juד�j�y�+'��乗�l���%��Q�Uj�$?.�����b%��`�b�؍�9���M�CH�����s��g�?�Mz�5��?�cǺc&���V��q�}�+�����䀭k�ۿ=al��G�Ē��ypC�W�o�������:r�-F���r���~V]�5��������J?���Y s�L�X:��I��������#D�@��s:���#���ƻ|��[7�����8���TvRS7�����b9S��lH;W0�}X�f�Ɗ���,nC:L�rքCr��8���#oѫp���##Dm���5�5���\��	�@^z����6���ռ! )���g�w��]ꅯl�u[,�\<F���B n���	#>r��a�w����dy�W�.�/�%]Nm8�o��P{��7�I�<t4���7��x�č���3��3�\��jy<�	� �z��2AE���y�į�!'ޗ����/�p{IT+��� �HDd��}�`���ݤ�q��{ӈ���m	��!���[O:Y�>��J�ȷt��q��Q��>O�+p��݀ �F�li�7\v;� �y)O������y�!�k��]�/�:@�\������v�D�C�ܾC7}ΫyR�T8�O<l�˙�����B��UC:�E�ub���&LqF�������e�P�W�8_�"�L�e{�k��k��!�Ϙ�cR6��g׆�a�q�ʢ����p���hU�P�T?�ޫ�l)���_%�<�~M|A/�<e�!}���K�u�U4_૝��g�̢Y�b��}b$����LU��V5ĉ�H@҆� ����N�oC�n:b�Ay��rӖ��i�,���*1������0�M|Ʉ���i7un��v����ns^�(�CG��4��C�s3 ������}�������ay�M���=^/v
���j�'�Y¥���.�S�Ԧ�9@3�[
Ț+{je�a�8h���fr��N`�&�����&ؼd�D?���n9�&('--���'2C$�	Ǚ7㬂�o��8���}HԺ�uL̉׭���~��2�L�|+�-��$��Y�1[����([�;v�r��N�t5,s��=i��;ě�e�"~f�O^݃��K����w����!]`����T�����h�<涅(�t�����*�_c�Əֻƺ?k�H0����8�����݀P'w�f��C!RqF����# W�uQam��{����J�s���+}�f;ݛ+i8-��ç�<I(��r��	�9�>��@ɪ!JW�4[�������μ?�ٽTp��#l��߻	aų"�����~�$��ۤ��q~k�$"���Ei?����"b}
�(D�5B)wH�@�m��9��~H���dn~,}���<��պ�����'��t��C�2�0V��P��x����C���k/oq��<׻'z�vӰ��hA���U�R���j��R���I�� ��Z�U�Y��\Ȭ����hd<lh �3rT9G�p���1�,NX���LV�K�BsN�����0І�jZ��5,��-�Qf���I�d�K{�'�)wu�O������v�˛�'�q{0Y|���:S���y���Q �[/`���B���T�rqAy�GVj��r��g�i�l`�f-IG��i�:EE�`�`���t��e*�Vg<&P������qvvo[GV ��m�U=����?�ed$���� bL{��{	6ܷ�ֿ��YyAj��L`��{w����p�׏�G,n�ݡ�ja˻T��a0�n��w ��+`bSvfJ5�?W�2[_���`��<x�7�7�|����pu`��H�;�[�.�s�eQO��t0o������j9���3�=� �:$����Ч���=?��"'���҉k�u�G9��YU*V��(�}J1/ud%֋E����z��S��2�������I܀��J��aLu����U�dQ���'e	����i#a�(�,�+�[��.�iU�����?e�_�y�6٫e`�:}ʁ��D�2���$��'o���,A*(�i�?��sZ@�JMJ���<	�ً*�#���]F�`��0��(���[H�u�|��쾁�W�M])g����O�y�`���Ԛ�ܸ�P.��P��j`+��p�80����Hw���i��=���_aɒ�-�}#Y�ĳ�㳶�{#�͝^+)e�P#о��.�	�h1�s]��ft�@0�LG� ��T�J��Y���cJ�$s���-���⑑��-V)�go��ei�%)�߉ʐ�rR��6-q�#�A�$�\�u)��	�YJ'�/��-�B��`�>�똹a���	B3$M�$
���)�"=�<��۽a�K�@z]�m����eͶ&S-�E6����o<���� �A���`���jg#���I��pG-��3o�����g�I?ݦ%�o�$��A)����[(O��ڋ���Z9�K�/��n�7�A�8�)Y��(w/����-
�ۈ����j�u��0_?-�f�R�n���#���M�v�P��:� K0��qX$����7p*�p��Tݺ�5�w<'��mj̰�ϛ��5�������H&�8lg�]�N&�^ϦD�$N�T�)d�;��E�I+|�E�Ē�gz�ȫ��p.�)A%�}�����n��ȿreެ�jo����׷B�Z_��ܼ��;��%qH�q����� 	G�����Z�x�}�����|*i�p�x��&[�#��:m��;m��m`-w�����s��O�o�;�^�\oV>χ�[���T��R�����\S�\ǿXI��6x�R�� �82�jJ���A����LÌ��e�rl��i��n�'�z-m�^�G�W i_��+Տ�U���ZJL�07k�f��X(��/nz�Lfu��+^D�5�1�T�q����jd�G�_0p�3֙�f'���c�M>P͝N),o�Gf?*�&���L�󑴛��?_���N�0�aDP�ت
�%ԿU�G>�L��wT}Eh�fDp�ߢ<�^2Oř��w_�n�k��Z;|���dg�Y��Xz��!���v'�@)��Ë��٨>��Oމec�)�i��oe���\vЇ�]K�UMҙm�(r�>�_b�`-�qhH"Drd�� �4f�(8͍�m4�׃�2NT����SS�F�@�Y�2d�� �`�S�Z	M8L�z�1�T��y��[�y�z�&OV��~%!��Jd8�.�,� �w�V=jE���S��mI�S����h�)yr�1) ��b��C���^��3{�ʥ\� �LS��5a�Ӡ����=�<��<��Ժ(�0k{xz�-G���[��\�������c��2��q��I�d�m��"jQ� `&��c�$E~��N����O [�2D2�3X��Џ���#m?2v�Ƞ�������@4t�'T�{�/>����O�+��	��`a����!j��%V�K-?wmb��pB[UB�(�F1���U�e}!-��o�PR��$�;#��ȥo-D7��nqN��%���K��Q�V�'3i6`5?m\:�
�A�4hfJ g^��lq*Ş2�Jy���=����E�%L��`�h��q�G����'�M�lK��p�z��*n���7�,	��oh����*��F;�r�I��*�b���Kj�&�_��D�pJ�B���'��4MP��cQ�'
�8p�o���"8(#��\��<n�΀�����s(vV08:�����):(!���m&�ye���(�o�&%�D��ܳ�? ����ceJ�Pd.G��WO����g}ؾ�6����`�#b��-�H�FO0��:]�2�$D���R������G�8�w�2,16����ย�u�q�@�%M_��kD��$ )�A�R�A�򨨘�a�_���Z��
}�_������n�%u�߀x�b�}�������W �[鎨�/m��V��Z'͞��ܤ('�.a`rdN�Z��k���q�a�x"T���^�7�Ƽ�:����̻����֪N�ɐ�hM8��?^�~�<A'�柬0+>�����~qJ-زc����S�x@�>�ƺ:�5w�;��/tN�%G��yŊr׃��*�O��3=q�$1>;��<�'�֦���c	x�'c��O�tĽLxR�n߷p��DLc�B*�׏�ί6]���$��?Cy��G��>�M9��'�k`u�	-"��H�������׵��>�"��ׅ���s8m��d�`���q:dM<�hY�\�D�1��C���Ć�&"�T-Z�%�� 4��i)@�2s�ʵQQa�C-G�3���O�R��d�t��$�+k� I�ڹ&�h?�����m�hZtLs��+��Ț�+�מ���w�(r�d�}�*&g�2�,S�A�-b�7-E���I.i�4{W�B�N�X�or��Bk3�NC.Q�s^,�@#9��j��i�Y���=��qqu���<)��h̿�LB�ek����qE`M=D�p��i$�7����-�|Cj=_nN�5G�����y��<��0��/���6��ܰ�Ny��G��
�:��<����JVEU���G,'U��YL�j�Eg�� p?�k)���[��@WK`�:�E{,E��dkLѽ�-��y@Y�.��J'��W������(�7����ԣ������u%y8Q=�7Ǫ4�k���q�d��w�zt�N���'� ��ܒ-C��T��Kk��w@��˲Q�����aEa}����-��U��i"�@]��Mqw���`-`>#��]/ҳV��ˊ5
N	�ƿ���]�w�GI�u���ic���&CT����Upx�YY����i�D��Յ϶D�7�K>2���&0Mw�4�i������	Y���""�V^S���ܥ��c�%�i $$����լi�������1kE�������x��h�M!=Os`���"'#8dgu��g<A�k�1�{�6{E܏;�1+a�,�98��rű���5��,θ�˗�I3�=�9;H��U;�}u���!�Yi�j��@ `E�;P$�[9��3<��f�5��Q��!lif�Oh��ȣ��b���6 ��}�k���ƣ�R��13������e*9��
�_����~Ɂp0��b��z`�W;Kh�4j�0D˄��B=Ct�",5��?�y�diK���B��ԥX�/$�**>�S�e��'6�ѳ��2��=6ަ���d��zd?̎�Eޜՙy�5q�T7A�u=}��]�F�Z8�5iB2AB*z��fH��*j�?��3E��=Fe�!��Ԣ%A�!�lX9�[ld�:���Z��yw	��ww	~��$�\_aC��½�\[%4p@9��;���W�:pHnT��P�E�>䂯����[2��KĠ�Ü�<� Q�����5[sȕA�u�3b�Pam#�UR�=2s?*���r�Ha����nsӷ��ϛ{��!œj�r�.T2Y�lݺr�D����-�أ�x�^,w@��Վf��܌"rܚ�f�B���S���Ox��,��ո�R�"ʊ��4]8�WՃ/Q�	WoH�
S��QЇ��	��:mPA����Ȧ��ɖi��Z��x�p¾��N�t�5��^��;$����!��+`L����`H�;% ��������K�F�H�Ʉ�1W��/�Q7�J��:s��!��n�Z]a��u�tAR�"�1�{?���d_����@x9��R*��lr`hX���Q�̗mlP{'�l>�3 �G��T(�)��w,l�;<����E`W�\ެ�2�"��V�u����?�h�����=��y��)�f/���y�wy[����?��[2A7UX ͇��4cS[�^��c��{��lwO�0�VR3�UG��U+�M:�GJ��ޫ� %n�F:q��йĝ�l��x���l��%���ʫ�Kd�>��>r�p�I�>��JIpsD�g6���иOe"_�P�AWMa^?�Q-��Q�l���8 �ͱEoD���d@�����%\�ϲ8�Vh�	�Y�6�[�c�p�����qty��p�K\f���Xg��W 9=׻�"��KR)1b'�6�wمsg�o?j�<x�9� j�[��q!x0�afZ&�wz���5�hc4	a♁`VT�<����_�����ԓ�:�̃*PM��Ý�V�zR�fol- �I�At(�Y.���5���`�@�����Z1m����ЁS%��V���m�7IP��F��6��ӹTQ�̘`
���k�t��N�k 6
ψp���ogj�?5k?��40� �v�M�&l�Q/�s��9�Y�tpe>Ǡ4S4��R�'Y�JC��ՂF�m����z�@���ݷ��,�f���:~@c?I�5�Eʁ���U�[�������ي����U�)�����$�KB�*�q>���2����0�Q��F�A�a�A��:�5ߜv�N,	0���Ge�<�i�����`�r?��\�r�6�I�F���O�����U�[�hƼN-aBc�(r��<j�=e&:㬀�5^+Q��9(��@S�F�����|�����SP�@UE��E�[h���[{@ �]�Ť���Q�����l�>6t7꠷���Z�?�����ܹOOYb�<�V;�fP�׈55���6B,,��aU�Qm��F	�����Ez1S���\�o�jp&�ߺ@N�S���{6dK&�=s�)<�}F�]�ĥ$1���A�%>c}wH�ϲ�վ GJz���Ԛ�Jp��Q�c!��XP����7�����Y�Y/\�\��>�ۮ��(��H�_D� �F��Q�)U���a�-ϑ�����-�]���+���䵧> �H�ԫjk��&�W4έ��vzRJ�n��W���q��o?�j�V� 7qy4��l>́ni�Фr3�F�W�n>*N_����m߉�[*����D�ہ�2]��u35����ug,�N���E��؟�L9X����P���*��2�X����װ���BW���h��-l�b�z����/z��I�h�%��w�=o`I�4ZCZ���g�UL�I1M�, ��O�	��0��li	��$�@%��</��7�8ѻ��r�_H��y�܄ΕQ�jVr��fOZ�*�A��7�]�����!�yC/-�5�?y�S/!P�^��hJ��S���!�A��m �5r$���c$�bg�]i�%Ͽ�ބ����%;��Nz������������ۧ�z���R`�*�e���I(�@��/�!w��-U���NZ��C�l]�OM�s,�����Hb_�D�_���p<� n)�Xa��Y�۪��d�y��7ץT�^��i܈�"fqR�~�	GW(w6m��V����y	��A�$��҇�����L>4H��8J�P�w%������I[����_�p]1N��PP@�8�Sr�(���{s΄��Ns�V`F�>Qu%Ɯ>��e�zg]ꃭ���Q�����q�|��B�J�u�T���;�ݵ�5*\�Q��!����):��i�f��q�� -�zE�ȎҴ\0)3;��L���<�@��Q��S��][��P/-�~Յ�rQ����r�eDˈ����Rv��O��8f�dvw�R����p�;.ѓ9oC��JҌ1p&0h�g��`�~��l�d�p`+P�[dT��R ��}�Ĭ?��-k�Q{CI�1m O�hp��-Q]�H�K�NxR2�3�6��l��ʨC��=gU�5?�|���3~A@�$s�|�{%5��9�"	�+D�	�z�L�C��v��H(�|7�a�c��\k�m�{N� �����萤�ګu'��;]�ؤ�@H���4��C&l%�8$7D�P`�oTw?���b��(|6�ml���B�S��H���`������$`�j�4VXU����QN�ؚ�gw��׳�_���zQ�|,8u�|<|�l.-{rA7
<H���	]��]k��}�֚%i8���@&�r��q7?$�C�
�m8���,!������l��c�� *9K1��g,�ۗ^�R�ص~�q�T�����u7M��}h�����3� ��.�r6ƄU��֦�Q�nO�/V3MfU�EG�wB-:�FŻ�r"�[�F�i������C�q^10�L:�Jy3�ֳ!�����H����V� �����b3�+�A��؂
����1y,?,��J��5Z:Q�y{ֿ6�6^j޹C���Ʃw܉ު���
߫��Q*���Rb�ͱ���at�vPJ{���Jea��^�A��\��*��H�`��(�q@[�,�0��o�3p�mHܙ�� ]�}Ø�2�Liڌ�P���p�^0y����d�&�;�i�/��`DY/�h��lg���P��lN�6�.^�'q�eJR8�T��$�#�87�f���7���cS�
5�Y�f��Xؒ@��v���uU��ձ�.�g-��y��U��pi��"#3a'=�aY�E�/�r�W����Ej�u�%q�O$���!-�(�ɒ[�ﳈ5nd�1��nu-�R��s�GON���LS�$WTfY�+��PN�W=�D�YH�ycW��ϥ-����w��@�ߌ���{̰��{��{��^e@�7�d�$���7N��;�nM�٪-R��3J�mH71�2�٫��+M����1? `�!ò���㥙���ǧ��I>�˰,����RS���&M$c{?�h�1U^��="��N4�'���ť��ޟ�E"�a莬��%nQ2���_��$H\B]qa'j�0R,Ia*��<����1�(�¶�po�:N_� ���0�N�AT"��U�%����ӯȷ��O�Tը2�}@�B*�7��A��aj�Lo�S����HUS�JH�>��;%v|�$��m�آ��}�h}�������x�[$���P���jE��xt�л�(^}���$UɅ�Rw������P�M�d>-&�FS)ҭ�s��m�S�rLG�,��3�/��s�����O�N����c$PO0w��N�r�h%�m|�{���^���� qR��`�L{͏;���? q���y���M�������m%Ø~I��`���Z	<�����P�1���W�������ή/�xN�Q$�:z��d,-%zg��H�3��1��dv;d�f<�F���=Y���-�޿\���Ŵ`Zh|��e��Sw���\h�Lᾗ��[�����u���I}�iX�s`�`'aS|ɼq��`A�Hc	� m"�ռ!d���;tW=>"�pB
'N��Z�H�7�
�[���S �������Y�k���ҙH���#?�Dn��a�]��i۠��JM�t3�*T�GoU�k)��F��n��sh��b(G@J��Aq7`�a����!_�;�����x�Pgد��Ô�/)wTB�㨽��{h�3��$Rхk�ӧ���I-4��,�Uѡ�;rj]�4∍ �&(������DQ�ğ ���G*I^{�H��2.6�-u�`���D���������耋��e_[p�]��)��>)֑���ϯP��G
l�8���h�J߆+0��ܮ{�4;���2 ����H�2��_�sB�<s?%8�6����ߗ�a>eD(s�3�n�m5�o��AR�_��q�<���hI�P��2\qV�|��Lx�B���t\4�M�;���B�3�T�����3��L;��jp���m�vٿN�}L��`궫奇���ea�m���+�m��y�sV��Uh�Dq�'��N���@e�Л`NH��Q���W	�<�>?x�6��)f�
8OScu�O�����9�@:���6d)�Ъ*K���s9��ͱ�g�U�5�3��!z�S���zD��.�S�����\�	�5��v4c,���}N-�6!s� ⸄(��S��k������WQk"#�[�D���\o�}Emq��u����)���|��A ��@Zݺ{cm�V0����x�e$H���+R�+���@�bgi�Y�{���sN���~��:/��6�$�Mzt`�K���D�o�I����S�K�8��E^DO�0��%���цykt�,8��nt�'�VjQ������Wd�.�R���ZF,���{f>��ߋ]SY��e�w�*Rߜ��(�jT���W�yaܓv�azS��ZxS;�u0���Wg�����M.��@j�n�~�'����A���,���o�܉ʿuj]Nc�:Z{k�<�����.��y�<(0*�Z�O��K]��{F���0����e��g�����f-+E���d`3�B���yէ�x ៴Y��CDa�am���υ� JEs�5����;���ɓ>vQ?WU~]cE8S�6n��T��\f)ɂp���3$B�[�h\zh����WL�����tro��v�e�hC�T�P�
��Gz٦��J����1�RA��~�2gk�a��!tt&��ἲ���g�⃂K�n�g�v3Μ���fuz�r�63���7�)Oѥ�-ea�Z���y+�T�����S��]���V6|%4���^����17���{*X���: E�`��SR$�S�(�ى��y��q�+܆��lF���@�7����+��u`{�Fzw�V�O
���b��2��@��a2�*NːS_j��"�pݻ�R::~�p�W�|�d�U��-9�W�1,�V�)��h����!ܮW=�+�x�:0em���̈́�H?F9��H�l�$��O^�.I�<7�Xo�b{�B,�0��X����k�*�� .Y� ū1V%�����~zKc��H��&6�/Q�=�HG;�>�θ(�Դ<%)ٶB���'���2��=�		Q����|6b��p7`h�|>s5vsz�8�f���i��*nb�U��=GޤqH�I�PZI��[�t�r+?[oU���5t��[d�s7T|��*�!r(��RZf���Z�f$Sf�*���?R54i&?�8-��/�+Q�F��h���;'�-eV$�M����ˌ>�	g���b�*�g1!�ԽK�3�H�/���-�!�~9��kC��ۺb�^M0"��؛BЊ�ļB<!`j�Y$����F=�y};�4�s�S�"�s�ɸh��O�S�S?n�53ϙ������۴��J5��f1�c,Tb�Fh��r��#p)XL���l���wW��p�~G��&���wx~��cA�`�U��� �����lS��<����(1G#�X1�I�����N4�t�Ĩ5�uG9�]eI,���\�V��^lK1�����r%�G��7?՚j����~���(Q�yM����µ����Y��c�j�Y�\V�h<�� ezPv0����8h�+1�Rw){ 3(woS/ڑ#`yW�#��|�����[f��2��a��	Urh+�k,W~�d��g}?b�7{���R�,7�U��K��@_C��x�[��W�˪A�jX�'[[���u�l�ک#Eᡓ�v����<do3��O��@;��k	~��/kw�\s�_����e�C�Lߐ�ev�O8z.�5�W?������5��>��&�"Gu?{��U�IKBC�)/zh80e�r�#���	+6��,�J[����n���!�O\:�J� !���V��Ɛ�.'�\Kс�z�_eN�>��⟲����;A9�HcY0��aU��<�N\�+(�#�!w3OW�B�8_Ҽ��^(KC���1� �&�F\+��=�,x�Ͻ�S�e����X�g���@+̊B�'u�9�w���F�X�P?����x�b)
QzZ�q~d�ޞ`����d�����{2�C�)1�w��w_�+��C����;~��Ɇ��ٛ��q���-�9��|s��J`��)5QD�_�Q��Qb7�d���a�@"_�|�&�����z�z4A��&a�>k}��9�C*+�`�w>/R+?I�my�S��B4��jķ�����f0���zi7z�s��Z��?��fD���dI�`0��7�X�7�����D��eu#��l�?������j.�k�5����h��(�2 �KgǤ���H@s�g�����ީm�i�+b��M�]�%[<�y�p�%�a�.bã�C�m��q�t�c`��i��AŤ����GI�a�L���%�hiYَj��J~Lwu�D������6y�����O�e�{9��I�z���Oe���� 4%�>�A�[�To��
�����O��X��Xe	-b��,=K޸Vld*0��^&M�xģ�c�R6��W���P����j0� f�|~����Ƴ{-��� (^mz�<��@����Tv�dW�%��[�����=/;W�axD����(ta�;�����,W�YG��
�	��_}���&��b:{,���f@P�?:���c(�kȱqa�sh�v��'��D�����Kt�x� ��R�
��C��I�q�>��/�����E��õ���'�j�R��`�x��|U��^�7T��o��&�9D7�W����"u��Plhw�M���� ���=h�:@͎1%�W��̉ի���,�I��8���5[�du�.?�}4��M /5fN�no�c�:�Qf���=��N�p Τ����1I�y����&r�ߘU�ր