��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ��%�͉֭�;��B����&Ȅ�xe=�ɫ�Y���(�A����Pt��x˷�Y����I�~�)��=�v�ˀp��0U�� ���b�<���
Eb�P�(�(=[[wQ�b���?�b0���>^s��m���4~������(����._[sM�Ғֲ�t�w KAL��=v��AP�b)�T��B�M=橐��[:��y�f�����+��-��H�B#9������Z
����5-��Kb�8�@� ��F��(f�un]K̀��@rx��H���m�	�� ��V����-�dȹ�f�
����֚a1z}�6�ltQ��t�������|���D�z�?�q�Ӑ�]�D��	���9G��@0��Gy�u�}��y�p.��;�J�9@�ʡ���4�9���@t�BܸX_�kʴ�5�\2q���!�Z� j=Zq��|���53xm
(�3�)+�����Iu����޵0��g^m4�6�Q�/���Я#ΰ�֞E���r�b*xۣU��T?��o�eo>�&wͤ>����� ���Lc��|6�<$f
���O�����y��*��L�����"/Y��iv�X�@��y���2�;�X�I��#ͥ��ӭ��&�:�����X t�4z?ٷ��X���q��1�]�V��/"G�#��k�(��v="v�K�].]d'�.
D��B�1��|_�D�j������p,|�k��eHҽu��M���x� nb�ו{��:L^�I������P�Z�"E(P��N���e�����4�$�0�O,Z*�>)Iݷ��:�v�z!Ϡ�P3����z��D����~��Eq4���>��wv�-�3�e��c^bc����]��J�݌P�������깢�!~��9{e�J>Bj�x	�FĽPSW�/4�.h{��]��Ì.K·�$/�E�*�'7���D�q-���Kb�B�TG��2{��_vO�B�X��Pc����j��͖BH�s<����Z.�Vy���N���Č.�4��(�ջ=�N�/�Y��k��K�BJ��i�:�-��]s�$�q5�X1��KM��/�ZeE&�X/����=3�/O������c��c��I�ģX�?7ۢ��t��\ym���ኦ�3�Q�!Z\��L�P�.��J�Buk�&Iyjf2!��w��!峞�iS�vQ���D�ρ���rOyS��!7�:`�<\��� R6<�>L��L0�I��n�9 �
������)��m��c�pU���k^@�$J5��D�W�M�޹V�tw��. Tv���wF�tT�!(ヮ�ίD6��O�;$ٕ�ؠQ��
����<֒_��SMH>�F��a	�$��|`ư�8�8�/>C�3��~��	ʕ&�ȸ�� +K�Ϲ���n���y�gU�Xf��xq�8E;	9�d�5��m��#d띅���+U�a�f���Q�[|ޒ�
�R+h��~d���
��R�k�C���*��b���6�����\�N<�b%|)gP3�^�#��3����W�Hx-��#y&W,�e����	��l{�(�K���?N�W�)<ݢ���m.F/�Ķ�ȅ��j�p�<>��cp�����=IE9;ޭ�yV�z{t
2�إ�f��*�� B���79��&�Z	���C�׀h!���GVF�^�>_9d��l�装����sк�s5pS=J��E�=W�)0\�Ďdl:�e��A�do�:[v�N~�v6��hs����"��� q�m�x��屑�d�J>w��xa:G��Y+�#�0�UzO{M��i���bl����8�����&2Gg�s�y?jQXHK��!v����+\'�_�'ǎ��0�K�ª��Xe"j.�S$��"vכJ�� ����s|�j���p�x^�
�D�x�*����xKjU�.%<t� I�}@���\ǡ{N�ީ��*g����g*�r0��� z�>�s��/9]����U�]�]F_�����1
���ix�F,[b�l�� ��X�O�c�9�S|^Kp �Ә�1=��(t��ܝ⼙��k��=�q�R�;�6Gr��^^�|�&\�[bBxC�g��}�K3��簗���BdF��ZJ1�o$YXlr�S~���}����� P�X���)�sޓ��G5��vM����G�{:�u�G���h��>Ł�Vg<3������!B�{{-~��R���p&f��P�="q����8j$�*�1 |Ά������N�cA�kH!�豘)�5&Nm$j��ɑ_�G�2��P�'3����t1�23�w�-'~Xb��u��pK=��6A {he��(�
�b�r .G�"I�?V��;b�A<7؏�w�m�)U!?=�t��[Ǆ�-o7]�p�>u�K�hT*B�(I��x�F���BJ���������JϚ��ҵ�R}Z��L �*��4��M�s��k�@���"f���<kZ�{$Ac���x����@��DO�ZQW_�(U��7�c'�0#@��'�Sw���vNS�S{�����9g6��
yplW���6�x��v�Dd6Gw�z��S�2|���.�AV[�b/��*����Qklg�Z��ԑ��Gk?�l0� o?�H~qLV��A�Jw?�C�B�e��w`cG��0ϵ��� ��|D
�ʂ�����Q�E�SE�B=�E ���_^�u��w�A�$���W[4�RRy���ɳ��t@��Ĭ�W�R�4�6<9s>v�}���[։��×�$N��x;}H�u�௚���B�[�$ �H:iP>��$�eZ�z�,�Q���&TD�(@��t������G���m����I�5� �y8:�#9�h���ۜ2���л�,�x��-�#�d�8��n��L��$%]/�D�p-���R��3�7W��*�Fj
���D'��v5�L<�|�lp��J�\	񸈑�}�W��&!-�b��K�i*���F����9]BuE�c���3!��h�|���=�/�Cd�Pn��ƚTߪ➙�l�_���ކ^��Fe� �y�06��ڕ4B9�H�?��}L��N��jC���'LZrO�5�"e�3�)h�~��P��WA%9қ$Gc�}����#�Գܥ�̰��uZ�0y/��!�:^�24�]ѐH��w[DXb��|�#~h �G�������&p�п�г��Y�"�(�����j.��!$�H�߱�?�F*rk�s2��3����bhԒ1��K�G���4U�-!/"ҧĀ�Y��+{rf�h���K%��V?�.��/w�=&�|���"o9�X��y�����DD4(� pV5�U��A|�1�t�GF�P�?��(=�\�p;���!r��;]d�����_���꒖B��׌A	���3<�Eح���8{��ʛ����
Au��A����iKmR�)�MD�*K��l��<)�]I�R���^h���>L�8���A����}�G�@�5�wY�M�kϥ��:�=#'�RK���iG�����ɂ��f��ӓ�Y Z;���3�{��uO�v@I��+ε�0D/"�:�i>��g�Uj�)�W/��	�kB����?EDJ$]���[p`�L� �0�%a��ge���Tڥ$O��N�����A�6�9$m��S�hF�8��h�"^�c�4mw�B�F��"3+*�4���/�T�u�C@�u�?'���l<l�p��e&u�'��a�1�e_���]-��χD�|i��5ѽ���\	�z��>�X�M	�W��bH�h(6�<��g�Ynڰ%M��%F��4/�`Z�F��P���v��:�y��T=��f����9/g�y�4Ul���c�s�C��3�1��+-;�a_�������]�U@�C*���항)�fp銵�:M��,���@�	m����V��r�P���SB#h���eA��:K�]�'�*�͐�-�M��`	P%s�����:�5L��L�_!*�9V����J�r�88'Ɵ���ʸT�5��=f�T�j�z	�"�wA�C���c�"��mV�Ѱr�g.'ܪ̓���(\]�]�X`z���4��Y�l8�tL0O7_�m���c3��D�ȝ����&���_��U�"W���U�oBz��5 =�A��D�!����/�0�w�}�8a��8�� I�A�Rq�Y��_NR��b.����}�!�(BQ(&�#�q��E)̲��I�H������ �D4შY.m$|��I�J�u�6��9v{�\qlD9��p�%��r7F��5W�"SBs�zf�e�P�g �L�iru�c �j�I��`�''_0[�@
�hf���m�3��B{�Q�a.X,WW���9��z�/�Qa�M�PZi��L\F�F�.��]����i:Y1Ǽ-)�����_���s�gdO]����\�_�^���VQ�z?�Y�.B(ׅ������m_��A��J �A5��q�q���q.2�:���m�o�g%<}��=�a闻J;*"�f�$|I�u��:�

��Zi�g�տ�^�+��P�.���3e�d�d*�Pz�y��o��)�<ډ�q�R�Z��(��o3?�:1��w~m��t}OS�m��ҙKm�NWi;�+ʞ;�����E�w�;=��}e�J�����pۓ�4畹���<���:�����nh^�=��紹;���R�4\�'�v�s?�� u"L�%l��W�t���r�o$d��̠%�wfvoh�N�Q+�ɶ��>���¹3VCZ}��F�&����8	�I d$�Ʉ.����ݘ�nW�j�B���Mq�,���Mj�sg�<x2{�7]�ފk�ф�����S8o���A�Rߖ���Q���jA����r��6Ҷ����K�d�A�N�--&���0D|�c��mY�$��#��4F�Eѝ:���f�k�m&lJ�hW�����x<?��h٘�S��s��C��i$$_�?B��A��+����"�3�{Cv�M�E�T���7���Fb�#���m�s��at9�C�}VƁ���:8j�2�����.GJP0�$�M��v���)�A���*�}x��]�$!oE�J�g��0V[�(��� ����{]| �r`P�ȵ���$�:r^�i��������;.��m�|"�.@]������P��&lg�)po��b��3���F��A��N�pi��e�M��<�����p�Lh�G��Pl:�jO�;�t��]:",����3�	�(�^��6(A�k?��i��V��J�wD�� �s)\����H���B)���ɺ�RXij.�[�ݦF̞)>�q��b�BԨ�&��[ׅ�+�ݭ�Vd�n��{)L���Ŧ�>�w?@a��_,I��۬�,�4���*S�ko�;_��oRfx�r�)�L���G������}��w����J�b"@P�O�� ��X�?3җts[#m�~�À}��#,�A��@�8��"�w�W}G�YY@ϰ����y�4�����O�Ѝ�U��̜a�K�h�)��1�e���?�δ镒}y�Y�i�[��DK}�����#�ĆLhn]�som���E��}$����(��W�Һpl�ah��?�q� �L��Pv��зi{ [&��݈A��v�?��� X���K��#����:ͷ=X�_9��YE%��Zg����u?�������B�2sEϿ��L�����H7'�$�`�������
�d|�	����~Qc�оx��6e��>|:���uJ��n;K&��ǵ7'��O�����א29�+D]��t�=`7~uk����=����[yY��E��x�,�T�~�����DY�r�,�G���FL��>��O��'>��R݌}zdl�Đ�E8Ȫ��@VZt����3���I��H��ڭ���6ı`��P2�W|�::/9��RT&��`�������GME���J�E2f!Բs7&��,�t��<�yi�8��A 2F��u��}.�Ri�s�c�*O�	z��4D���uvW������Ux ��{��/��:jE��~��T��8�n�:}��?Swą�]�2:|R줍npǥ��5�ee�n��pbڇ��O�Q��c�V�u�t�		�Z�&˯�����0".�Z�W������OƯ��~�8V����>��*�g��.�R�6�c��#�����!# �;�{�ZN�l��Vo�B�X��\�m�ѫ=ith�{eUR�u�'����S�ʧ@u��n ��폊�/Ʀ�瓘�{b58����Op#?ow��F�T��Cm��Í��菂B��or�g�_Q����X��=�ߕ���ʭ�X� Y�#�&�u?��~������sM�S!3�Rv+�!�M=��p��?������c�1o�yyhY�l������q��.�̹5b�� ���o��B�H��_��rn���!q;�|c2�d!�X-��9�\�.�f�
�iZ4�����[@�$繫�'��(؜�4��zwi����	N�������V����ΐ�U
d�Iz�q=h�3���R$�^bV�yY�'�����B�0��[3�+��H�������)��b�+_�Nf~W��]��eͪ*�Q�'�
�0�0t6�*������-�\2������:R8w^�H�����A����+����%�$�n�*���?�����D�/�sR��wv��f�D�k����o�g>Q�!3ß���֌^��5@O�!ߓ�������S�4�4E�J�4~Lp�^u�:`u�E3�-li.��L퍻>��	� ����of��6?a�ߦK~W���5�b4����b��T鐾����t"4�8q-I+���A.��s���u)�M���\�"d��K�U?�#��Fuj��aUpłjQ�5HO�ݫs<\�gLe��|7	���j���]�­�S\��mqg��!�������ޔ����� ���LrZ�­�F��`RN�۠�MҸ#]v-��S2��Q��G�������P�M9w��k�K��?�#�\\5����!H��j{�`=���������-q�܄���"^]��S��p1�*�bcE�����_kz��;>�k$"˅����@��&(��? 8��[j��8Rr�c&9�rp�P���$�s��m��ߺ�3��E�E�g  D������ 4#Xҹ	�	ȹ;��
���9��3�+�^�d���QpJΔE;�AeK`"�w�U�o� �r %7H��
+v`�jT@�xL0���Vp�6����	}�ICc��90�a�g}*�,9-Xp��r�?�08[1dyx؅Z��@V[��2Lb�86�Q��E�U'Y��)ډ�N�q�l��Q_�!ዀ{&ƨ�q� Ĥᰇn��2?�����[q�l�b*Q�^�/����"�b��f��^*E�⹐WA�;�.�I��e��X���$A�\�X`w�:�pD��6��}r�Cߥ^8W�l�|3��;i���;k�n���"�	b-*��hr�b���
�L��A`�,���/.ڑ|��5���2�6�b�AT�Խ�g<$��|��y�������,�RA�11b��D�p̗��[��2�F+I�ղoq���p.��\�"��J%,��0jAV&rb�e��?'V�t7�Hd��4���q	" ��"�HT��f���`�XG>7s���Pg[�J1,^�B5��_����''M�������7���� �+��oץ�a
��B������W������:��Z�0�{G"�2^�Uz9�d���E�ÌT/���O���8>u��2���S�c�6�j��B�V<}u��,e7�6vQj�1�x�ZJ�M�B%_~Y',E����@Y:
8��B%N�΁.�-І@��"���b�@�T�F��	�����r2k���|]�0%̅g��ihP�B8c�D�������Q����L*�h�Þ��=�G `D���@��/�g�k�b�TE��BJ�3me-.�ԇ�}�4�a3��<�E|�GIǣ�7ł�r@� �FW�-¯Q�?�O;���Kj7�Z�P���P�X�<�e�]=��;�Ϡ��}�j��kSv_0f���dZ�"����E/A��O胛s��I��Yh�PgEC@�=�JܨQ�,P����B�I؍�,ڗ�Yٯ �О�r��/E@{]��O�P}x���WqD�r��B.�9��T��i7��6,�����K��6�N��V����YGc�GȌ�Ð�����Bj4w���U��{Ӂ<�t:��+T�Dwb�ѕ�5�k�[��Q�q.#�M� �*a���J��K��fJ́禂����Uק�4Qzk_E?��1�����Q��U��,�"'�r���W�� M�g�z��rh�k�Beш��OqĀ4e��~�f�Q�lT�*��ʟ&,�[dL�>X�<د�m��ϯ�߂H?CxU���=�9��~P��w4}E���-h�
�������j����FJg�ڮ�褢�L5�󤸵���Z/k��� 3B��ܲ��qU��D8ʹĬ�������e�8�=�99Kf쟻�y7t���P��x�r�FĨ�8@0��nه�/LYr����M���u���P�nS����Q���4�Y�{�����w�#M_j�e � �}KWp_��1�6ߏF����NΘ\w"�L��T���h�v�h�P7��[��N�ͳ��"r����l�C�=�<����G��vUŃ9�y��f�� Zwu�҃��U���<���0`���)�bfM%w�dg���ZW���3'22�t3lS�b��V����ч�$��;�롑�{ ��>籕�p,|�I�hI��!��G�
Bc��].�j,���n����r(PYU�^�� k��B[k�0���1�`��k#��_T����_�Y�ͣ���Bj��ɩ��a�4�&a�2	�/�X�&\�V6�1�����N5�j��	�Z�	�;N�
Msn;��%���Ǥf]~ �{��%7k� �~�rj�VcI\�
��d��Y���iMB����֙�i�z��	HC� ��J^+'G'�,������=)X���8T,�;ʱ��n�M�o�7��TL��E�^�~q��,7�P�ʎ{�=�P3:�����d:�����{,�h��w�]����U��q���t=���iu��H|H��KâZ�Q�$Fm�V��t
sX+��	}B7��]�����B�8p;/4iD���p�L��Σ�r�a�-!�Þ�z�z�qՕ�C�
f��$fi��}�t%����3��A���u��FY�I-�`����lA*�Nt��?N.�z�\/���� �k�$H؛��]d���9��(�e�"a��+���*;��?r�Sy��8"�WM�;Q��ay�&�5͈�,ח�Ծ�;�w�S�L��|Ie�A�k����vdՕ�~_L~���o�f(�de~��6�`.�]�3�ab��_�A�f0އ
^�9���Jepݮ�7�S#��������3��\Ь����15��,2���+���5�I\l�(�S��6�����yߖ���V�-X$'y��G>��Q�^񯀧_�{�~[�/������(��#Z��5
!ˎ���/�p�[D�E���h�؉��&��mn�����+K�;����j�����C���r�9K%�>�Va"�p�m��qP*�T�]�!-F��N���m�.ed�[�}�]�@�:O���9�>�DN0���'f���k㴇&�[TBS���c���x��N��C]Ԩ���Upqw�`��
9D���� �Ld�,un��`�Y����ҡȽ�g���88Zp�=��[rliEEć�VDʌW����F����	&35�����2���Ǖ�xLҴ-����g��4���\w+��l��F>�P�BIFt�=�h�&�!�+>�$ g{JN��ꮪ���h,�GaQ���+.�+��Q����W��T�ʮ��R/�͉Ȫ��Ly޵E�JA8�s?�F�Ow�

�t#Ass�?��ʠ�5�4�oods�j��pm�/�}PsaiS"=����\�z��<g_/�p�=�g	s;{���u�����c�K4�ŝ�̷NG.ա��-����-}�b���d�f�4<䩁�^��F*Ʃ׿1;@sP�Y� c���QA^����Z~�ŊWk�'�%�*Wu����W^Z<�p�w��X啨�PH��y1����󁍦��2�l�M:��%g1��jM'ϐC��S<M|@�;3�&�$�Vֽ^w^#��6��Z3��q:I4塁܎�T-���*���S�=��_�KĈ��P�̦Dt�$��u��̬�7���E��H��y	*�b̺�G��䨟�'���w��n�5�"�-췕ȼ�n[�[qu����*.�ZY��=<����'�/���o
f|��߂?m���V:��I��?W0�Uy*�]�h��1^����a񪀢�0H$a�~q�甛�v��ҫ��١E	����s�����f1�i�8��"����R�텋��F��9�y	=;�.�L����G���\FE��&:���>B��r��1t�zz\��{:v�d?�Ƃ��O]�a���N>��=��֌����1q{�JC�E�U��,^���Tb�@.ViPej|a� 7�p�`By�TX+��-��>!�a�x��5����B��Љ���\pt�?Tu�?o0Ϻ��/��ZU�SETd锘���\BX;��������٣{��t/ۅ���Q�pL�N�fO����T�H��'�g"���`؞JyB�H����L>�+#Z����L�T�� =������`���'F�F�;A�r*�B8�^͕rTՒрx�c2fL��b/(���x	D���%�~��J	Bf�Y��C�K�3�}B��Z�i}��0{i○���4� �!E��K:�����O��s��)�]�H�j�~�K�������&Cz^ν>��C#7]�ֻsi�̲J���Р�U7L��ꇴ}��
��B��r��w3
e�9L�}�}���kq�ϔ�qa�슜�[_��������#۾�E��"ϋ?w@�9�(m��
�P��&n�]��MŇ�[�iq��k��������t��֌\䒗�!5l�\�9h�AG�g�Ed��ǰ��n�-���-�}K�S,(D[W>��ՀjSChN�9rm<W��o�T^(V| �h����ĬlNt�J�S)~k<�M.���[�i��VBk��h�V��àA�n|ͥ����&r('�= t�[���YD�ܲF�.GLh�43/����	thX�&�w���J1��.�/�nE��*ȄG������Yρ���	EY"�Vi7�C|�2����l�E���~��k�]�y�!&$u��u-Y�&������9V��U�p�I�����0fS>$�[w�+�K_�k����=��8�1'4!1"[�%�:p%����0 ���}��dN�>v��q��qo����4_�P�!G���{�&�n$����$��g�(P&��m�:�Q���@�*h��1n(1-�e���ܠZ&��)V���R�� ��~<���h�tg����/Z�Q��"Z�U�U�������u���]��hd������!De�, l�KH�$�oFj���k
:|S�6#!w��Zb����נ�%�H�fԌb��;�f�^j���]�dV�|�LP�� ���r��-�N&���@*�ь7@�D�Q�*��	J��^���B�ΉƠ�7�(��� ��т�4��:���ؽV�Q+�A�L�5a�U�9ߊoqox�Y�R"��)d8Q�������Ѹ�U?�
{S�j�h,��u��V�|)o��n�:���À'�M�A�����Ad]��Q2�x�A�[�"����1_��`�YS@�$��0g1,��\�&<��)� ��V��KF�1���:� �s�Q�"���Y�p'9�t�pz\���ћ���盺Ò�x�H̓�	��㯖��rA�Y���m�Ry4�ȼq�׫~�E���_n�F��/n��!8����d��F���\�0�z
�C��6^l��	v]�~֎s���K��{pBj��XbE{�I*$ct���_�T�4�eĭ��ɂ	��A�l��hW�,Qĳ��e��<n��KD�3��$Q�2[�=��q��{�$��uPV�����	B�7�)X2gh
	2=�����V�̜�fU:.��}m�5��t���#C+>�¬ԛ�:��!w+Ρƾ�\o�i��Ծgr��رvM�����u��d�����������8%ѩ�=���? #0�����ƫ���l[,�pK� ���V5��J�%QaF�@��Iʘg3��Է��y$�Cv�׹���7�ӆdn�Ȝ��q _,؀Su���y�ݲ��>FlA?o4`1����q�u��␣<�؉���׊�1�s<��BiƏ��'���^���ᥫg����n����Gd��Ph=NL^FJᅬ;��%��$��(��Z�v���2&-�(��X�dD����R��Y:�������LT��FRM>J7���TJ��]CD��dM�e�A��b������Φ)�&�v����yoK�'��p ����5�:�EmSo�P������A������7@�Pp�JV3M��{;R�\�+M
 ��uE��⃿�q|��"�I�|��ۥ���w؂��Ϙ:��a��SΉA�= �4�1B�.%i��J!���e4R~bh	Z�mR|)� Z{�r�m����1��Ex�ɊL똓&���5�0�/���N�0}�4&�Ễ�Y. ��9���iK���S�d�u�����6�uo)�ѳ�J��"R�{3�Dּ�z"A\� Ոy�:��(SY �|֗*��.1�k���T�WIB�ޯ��,���J\�R�1Hgf����K�U�?���JWͪ��(<�V�����f_9f����Z�CO&Q�)B������^|� ݏ2���v��Q N]8ftcP>��."L�q�h5���aAÏ?X���?��[�#�I��a�������$��f��x�bw�'7|=������2$��ؕo�hrÓg'�J��t{.�〗|�ޱ�� <F�D�����V�j�<�Pc�Bٰ���>�6����>���"z�����V�����"��|��VtV1����3�]�<�9\��Ȅ���rf����	��W�.��,ۘ%�����?)$�k��|5Pƈ]K`wY>�� [��@�pW}/%�Z�t��
�w��4�~l�{�	sGp#�.5����� mY�<K�A�l-8�b���7w\~�E�i<��	J,��5C��A�4�+�Vo�v���q��p�]�|��@��=��P����*�L��W������c����`{�Ą����m�L@��>��tX������0y$�&�2���j����nK��P�-\���5����IB��-G3��	��@c�����%��j���Uj���`��Y����)B���\�{��B{�['F���W�M��v$�k_���	�P@#������Xd@���SQ;�/��y��Y�ߞA�oE�T:��
%���#�/��($K8��H n�BX����n@T�[�����������*&eH��+m�qA��U�	Ȏ]��㭣Ѫo�J�h�7?���<F�߼�`#��A��{��L
�9�c����uD�� 8�W�P'��T��0jr ��S5?2>gIѧ���G��)^���jvp��B��j��9!�����|�F�R���ďc �%_&C䲰�lNK-5�_��I�y��/z����a)�-a����8]0'2BHj:��],��ɴm<�{��`����|��L�C8ф�K^%;�)��@��W�x��7�)���{� Dպ0��c��p��b�oXL[jN6k��瓅�2
�p��Bw3���s�V� �Si0F�f5c��cX�Ja�xR��2\{6ǆ���G&U?����	f��T�eU��Gm���+t%�%�S^��ǆ���
�dW���qF� fmW%C��0Jep.
av}�b��#��k*2ڪ�Sa`��6}ˑ��)�[�o��JƠE�S��nZv�W[�P�܇|�|k�p����K���g:y.�M��	�����:�c��w���S��Li^�8��5�{x?9s��~gD!i8,����]p�0��ʺB0���vN�]��ճbϣ��6���D]IO�k��Z�\]uҾۆ"�&Ȣ�\����DMfDakʴD�;��Y�
j$��k<������R�2%{���6��.y}���$6d'%n��˪#�����O�4��]n�P�T�SG��x#�K�:;�3��P�u�k����Bh���1�t������u�~bOF�Ԧ����,��˟ǻW����g0è�]���-�ܦ�/'%�ƽ����x�7��)g��u���O�(_ܐ�%aI�?6#�k���aB��H�6�\!��q��b�ρJ� ���z/W����Ӑ�-4�A$�.�.��B���5��.~�H��@��晟>��޺��R��Ho�D.>�sl�%��Df��LV�@��;Z$Bf�`��m�����AD2ɟ��Z�݌=z�]v���Y�%�������\,��m{=�Ss�����[�z����@䂠�`@�xBNx̉5t���z���G�����V Y(��t����jI��C��U��C��+W���E���*�Pqv����Ѩ�����-�Pkh�3���ۋ}{Wd��W��#�H�@&b\)��/���L��W�"�$�TV:U��>0��{]Ժ{�v��~��u�C/�"���7�""e��C�0jl�����EW��?����{S^�����k:j�{�$7�v��|nf�cؼ��������`�^ɚ�Z����_�����C�P��ډу�ӎ�Z�H(T)�)�{x�_x�B�0S2e?Tm����u~�R��3Y9�$TlݚJ�N�Ť��w���W2ڧs�"�ܗ�f��N,�]4Rg�֗�Q�h��y9�N��������x����6���:��|�Pq@DS-ܐ���b�Dm�p�� �OQM�������Z�����Q�_b�aK�K0W�l��ӱʬ�6�L���z��=�<9͙G�9}�Y._ײTy%P�VƎ��(���h׻�LxY��J<z���t����u<�{�z��{o�� @��\�q!~�I=��ߵkT1ܴ���*|ڱ���ys���m�1Q�iD N	]-��U]��?L�Aa�0X���
���_��#[?{f�9
��6��&��n�?�v;Eh�=�ko*ui��j�&:�=��&�Y�[���S��r����`=g�T�D�.�,o%ˣ�,6-�����f
�	����jW��l��0��,�w�T�<T�?�����D�T �E�E�B��n?]S�ۨΞƪ�����&�ť�&��[ <��[ߴ},n9x��óHqr�;|�K.���z	B��k˼ ��8�����9��Ў��h����,)�q�ͷ���\�$ł�J��ۓ�Yy脣F��^"moF��@+d�����cW�%�Db�R��Lv�x�=��՛�<L��:�a�}�U��Z6>�hH�I�;&��O%NTb���D}k���c쳯]y��Zu%����`���.�3�cCod�n�]��~>|��-�_�����E�[�̀��q�
�Ġ��h����ܾP��.�N#GL|��PF\-�S��� �)�m�(�<,N�� Z�m��A�R�)�&�����`�~>��3 +�܁	�6��&員�ލ���pw�+��\��k_A4Q�Z������n�vZ�-=���\��<b�J�' �B�Ӎ�>m&6*�.O���Hh��.��Y!M/�KL;���Y��B�DHE2���eg�b��-0��]w��b�G�mU&я	+�~��T�8!6�cBGU��h}CP
�"��>�9��F$@&P�*��'
���-�"��e*��)�T�Ͳm�s [�!0�E���7��AI����U�	I����:"�����?�T�YW<��|U��+�%RR/��u��U����W3c%���@�)&���[��ͱ�9C#%
�X�Z��{�/w1U��!�!d��MtI��zu�t��j�Q6l4'��U�ܩ#�!~k)׫9�Q���
)�75,6�&�_�� ���9��kzø���'�}u�Oť�\�J�z�1��섥-ǲ1�˪��.�G#'!Q�|� mf/7O�;�i�;�5\��KB������XS��l��/C�G�hv��i��2V ���am�4ҙ1����;��OB+�ZpK������h���wun9$����B�I�a�:[�Q����b�f 6�hT �"�7 K�G�{FVR0���V�|)���^n���IH��*�}�g��ޙ���ģ:�an�m�ۮ��Zj�A��t�#�?���a��np10}5&������$ko��Z^h�d�:W&�����c�Yf@OWC����ʴdu8f����"���;��0~�_g;h��
[�X ��a|�#3��������;�v��؅[o~k���N�*7�\����~��$�tnP��;$�����r��CA�[�ߐ��)e�o�������]���JX���N�m��BEzZ�P<KJ�yׅU�fKx�Gz3Ⱦ�<�`����!Q+�{m$�Sn����\���W���V��!Q*(d1���ũRل���� �KH8�æt�`���� �DKq�4z*=&M�7�2
M�K��!�]�T��-0Fhp�{u��4]!-m�YdK�p(���^��Ԭ����������P��tw'1�����[��
��8O�?6��BX>b����6$����e�c�|�#��LA��_���ȝ��<E��H���"� ����Vh�iٷ�8�AA��M��^���ߡ �Ya\���>�6����Ff8�d9W���� ˖4���Q�?�����m $��`�lB
�H�����Fm��cr"��p����Xb:Ѝ������`��e�~�6k�6�p�s+�y���6��.�k���������#<l1_-5|�S���x26ƦM�&=ET7�6��x�T�r�\=����Z��*�a��jx�~��}�lˡ�v��1��6���;Чqm�����_x� G�<[��Z�'����]Fx�'����!&Ǭ٥��yW=��ah��d4�snq��}��
{�(?g*���x̼�Ǹ�%D�Q-	��z!�MٞՋ��R�F�~��!S���m�"�-�P��B��K���	�s���K	�U�D�����ZBl4��A����?���ks�ȩ/B�0
��	 �$|�y&6�p���:�֏x�Y��jV�QX����fĽ_�?<3�~�B@����|���L��N�H`�޸v/�5C�9�Pq 8*��p��l��8�����}�M3�L�Ti�ڡ�LT��ӝS��qV��g��z���$,7ɺ�̔m��kl߬��~*{��~-��u�#6�ƁXVŶ�1O�W�=�P6�鞑�O���N�h��Iz}eZ��*�H��ܧ`������-2B4���q�}�����fO��T-�;,wC7�x)��� �7�i�5��B��GT�Wk���|K�����Rn��HI�'�!�.���i�Xo*�f��<0y�������U��2�0C�%>Ta����~��l��(0�������C�f�,ۛ���);O��\����R�i���8�M���ȳ��yK�IX!����TU�-������	 #����Ѐd=`~y�i%��	�cR<�r�d�:��(�AR�Y����y���3�-�T����^���~�l7yv�h���@˾m$f_��l�5�ph���g|߶Ϲ+�0T�k#9`��v�x����t��>�ߥ�F���y�0���W����	��e�̉՟����S��ȅ"\�5��Ny�d �@���A-i����d��1B2��o7�%�F/yG9^����\i�Z3[v%K,Nx�g�������w���FL=�@��f��u�j�_�K�������}�W��c��'�tC�T?Cn���]\��eN.�@A+���h���!�S{5�2���8o�uXl��v	�Cu�\�� %Mvc6	F/�Э���)!�æcy����+���z��X�J�ڤ�`�#T�`�	Z+�e'	Ttkp~!���4)Ҝ�X.?zYC�LJAMTy�R����fI��g���	ŭ�ʭ6��.� �O~�������F;e��I��f<��T�j�i6x�wr-.yJ��7ة��p��
-{].v�3G��~/������+�
u�;}DgO�*xmX);���qv�ΎH��ߔ�VH��=���_�@���A�ŝQj}e}x��qy�e�6���
�� D��N^J�1��j�NU��yx�gn�~x�:��{\X�0���EUcT��F7��S��G����f��涃SIʥ5���0I�$�
�]�b�4��P��xb��B�
������,�nD:k�l�R9z���6ʤ�o=�6�oF���㤣�*cOʽ�c\`��e�=2���3@<�����Le X�T�r$٥��STKN2k_�����P��RJ}��զ9 �R�ߛ��դjmJ�+��x���7�깤��@���g��b�ȭV����m��_Q�g<0�
���Ȕ�"�L�ϧL��1�3�c˛�SOwh�i�_(i|�ԌfܦN��D���YQ�y��ϱU�ȢO��3
Pog���|0��#LWdM2/�%f��~���h�4�(�o�A�:C���\�����Ub[���U;5?� 6�8��6���[-!]�̶d����kfxx�O+=���$��lm��X��ɉ�L�W^D�q�w+��ub���Q�QN\��W`� ڂ
��ɩ�M�L���0��eT��,��i�_7�����Jx��>�W��6���*�СL��Y�	�0��^�d6�X��,a�:����)t�����ՠ��������#�A�"��9~$�YA9���v4��:Fa\�#d��7��0$�*_�.�$�K��}�;P��5�G!UQ���s�}��x����8`���ע)h����'
�@u�:ϛl��񃉾�s���L����;wZ���,lp0�k�}�Đ���c����DEh�y<�&D�f��b�_y�T������,��S������1��!�^���ON_T��<'#�7+��L6�e՜��~(�8w��E2e��7�����;�$0�|��6��9'u���w��GLW� �˷nn��O��fE��¯
T1 ާ��U�\��\�߀0%p�8�*�
U�Q�k:	��Q�\+6�ܟ�],7Y�
Q�u��]PU��'�b�Ϥ�9G�W�G���_;���m�-��A�S,�`��CV-N�'õ�X����	�����?%{�!�K'c�W��U}u�'�t.Qd3/o~�A��1V���=�:	�#}�[�16�LRD@�L�g�#q����e�.��,�����Nc�E�.�nÜ�sqYkT�k�FO�y�/y�ޯ��'ߐ*��]�"�x?��@�b�ỳ�
o�/�$!��U�y�.���@7�.K�|):�e�/y��Į��!RAK�³�X쵯I"o6�hBXL{��,:)����
�W*�Z3H.{��E��;�5x�d45/���Ճ��as��	��){��5U�܁�j�gG�5[k��ʥj�v0E尷�K#��]"_?I��K�Q����U��+��;	s�n���Aa�i|n�����cwy7�_�e�Q����a~+'A���=xl��4�d�:9��X�y%�+�$�o�8�>��C�vp�@M����<<^��"f�[�g��l���2 N��2^f ��X�w�^AI�H�ԙ.0���2J&FAt���J�#�v-�U�z<u��h-�!����ˏ�T�a��3���lrؖ#�i<
ϡ�i&`̄}sI�2��i���M�r��Z�9N:+��F���s�s<��`>��m��KƓsSΰ�ߜ��s:^�����0wB"N��1ŵȉ�<5Uq}���z���\Nv;IP�Cn�G<P���
��A��	@C�Y�H*#3&S���`��#���pϾp�Bj�qa��>n����H�tߚw��V�Ow9""I�u���ZN���7p_�u�w�2�|���ɷ�Q�����mSD�V��<Q @P|�Op����3�5_�Hd����8��!FZI���G��Sh���M��33 �:Ui?oĺ����١MdU�Vy!Yk�A���h����_�~�m��h;������8��F%���vys_$��h�=G�^V ��X��-��T���~)j��T3I�9��eU�&�����Uʒ#���?Z�UL&��[l�8<�8��]X�ß�)�Z�10r@�P���Y:��+��6*����&P��G�Vi��Y���5�ڹ��g̅�:�cb>ׂlÚT{��u�v�݇~�!��?gOT!�#_�"�W}�\�8̅��ר�B��r���,a���6"�ˏS�:Go��"�=�24|�'A�v���,������K\V��J����VH���@(�6.��-�Ħd�q[���@�EAwUX�炰6��U4�a�#�J� öD�a������`�b��O�G�2�NЮ�i�XiT��l�_��K����	\G���H�L��B�j@�I��:�p�d;z|c����P?�3q�tC���x��S��(ڼ�v(\sV�b4��6Z�ݥ�o3 B�8ML)����[���5�?��';X�}̧����Y�+a��О\��|��f��9Ϧ�ί:CJc�_K}~�@^��k$�����O����Z�jF"���*����U�g��&��"�0��-î��Z+���Ǌ?���$Z�Vt�d!�n����	��R[�H'���Ol�;�C#��
Dhy;q�*��7�����SQG[�nx��>�ְK*g���n���li�9�Z�Kܷ�S�I��]��8���-DoS���G�p�*_!�S����*�A�V#$(��!8���.dR�f�?����k����`Y��Gĳ�/�N��Q��T7���߆k�8����h �H4	��b���Eo��@�V��;�v29��n��/�.|N��y�X�+�ȸO���!�
Y�R-�b	�hM<�;�`x��i�-��y}�Ј�*$xtQm�?0�FcNB��0k���Э-7�n8ǆXh�	S�Iz3y��nO�a����؞�r^�e�X>�3_ ���㺌#�ǎKb(�
}E/����#�o��'���xݐ��.����o�I� t��b��s��"��ٜ�����ß5QE
�fJ����������8��FΚ����ל��n�e��0��TOⰮÛa�k�}���/�ū�M~���T(��R��qE�)���XI�qD.	�$���!�'�^�7��nB%��0p��}M2p��Ta�����޺`�f(!WU����=՞����6#��r�?�?D��Ki@�n~ �d���C�k2Rd�e�ۥ�����(X� ������A;��*�Pu�ǡV3Kۡn��7Ap�k�<8& �5h!g�n��U�X�rܟ��YyT!bɨj�WQ�)�㐖D� �&OB������q�憨�:�6NvmyJh�������X��D	�ZW3~̈́¹��<}����#f oc������%��'�?9��!��4�� �ظk�"!4��-�i�Jz;��K[�~00C�L�]���a�*/ �	��w��J��g�����4؏��+ ~�=H�
��eD0j��L^&g��UB� �{3��ٖ���Jދ.Z��2+���ܰ��m��YC�{��#h%]7Z|�8�:��r��wr��e�����-�dSb2����޴���)�N�������)��gс��{�♔R�;���y�V�e�J��)Jv��Z�f6D�M����*������LW[�}2�
0��ԯ��u�*7����=67�۩S6�;�������=>Q���wLDn����7K���ݼ�����K����#�5����A(N���t;m�j��$�m&��`�.�Z>b���DD���Ư�YT6Ξk�QrW�%m������G������'ʩ�ᅁL�q��x���'H�
ڥ���%x���	�U��E�Z,(��eBșfױj[A�Gn[Yg�[��L��x�]1���� �`��=?��\�5y�N�����	�q[˱�V��4�o�������a�����\r
�3A�~Pj��E�5�[�q2\j�g��K&��c�O����c-׀р�5*�l߱_+��-7�A�7�����މd��;򸞃#����>=�XaG��=YIo�j[`_�}E�|�%k���z���-)ls��Rg�ζ��N��U	��,����Ɯ�� r���ٙ:�l�`�.��XlǛ/JA^�nqp6�4,zD�i�E�e�7�_Oo���2���
�r� LrqBQ����t�l� G=��Jy{��ʚ����]Q�jV�~'-�V۸M.#�)Q~���]o} ܴ8ӕl�O^{Cf;ͽ<�ڊ���O���^C)Tk~nhG�;��H�I�W�[_�#���Q�`���ѯ�K)�|Y$��Ū���kc�
;:�j*G���H��������-QXe]_6oa!?8=�O��]��!F'�Q��¸6a��l��t_�κ�])����OuY5�q���Y�1(W1R;����/>:�iTX�����<$������ܓ�hm��Z�q`H��WEG�6IH��_���wvF�>�Ս�����9�wX�lΈ�ACwȱ|c�	���M�ʩ�YH��ģ�F��a�$��|Gj�~����vt��%��;j]�4<���i.�H5M���%�֫�ׁ�u�W[",/9ڟ�/��,zf�5�`{w�  �ä<�
��������� �y|b��8;��
4L�
rr&�
k���F��.H��9�研�|��kwP#E[�܏�ru�lyG��h�֕�;�GY	�VHwKo�*�U����)�"��/A�
�@�+��ֳ.NY<�`�=4ԙn{}f(�j}�zi7k\�SmN'����q�~FQ��
؇��]�n<Qp���
�x�B�RB�&��"-��^��k�T��7|F%�;.��/����pEӫ5��y��۝&A��T.�C$�j�o|t���̣z	fgS�vL��w+���ݺ�RcU 5��<p�!^%�<Փ�4(�l-�Y�㪟8��R�P5ח�;n�w���z�̲~��l�6r(�LlȰ��I�ƴjd�h�7z��@K��5�L�ov?f"�L�S��� ,��*��oL<�z+�`!R�AIl����Q�W��k3�`���0K�ii2��o���c�d<�wn9��Č$4l�1Xk��'wiuK{2�uj��	�y�V<�ӯ� q���,n�T2�k���
��poidi�2N�t��ki6M�p��?�����Y�MP����D
���^%�pGB^�;�S'c����甙A����V/��;��m�˕F�DaAF�x�L��e�8PQ��:Ā�o�35��ԲO+�ԗU�
/b �(�����ʬ�!F��.n�y�	8�
.1�j�P��P/�u-G](�i�{��tx9'�d�RP�ԙk�W�����	`S�`�H�����>3�n��U�~nn��HH�D럹a��[�ǚb*e��h+��W���P��qI���0�ˆ�V���_.dCbdC�"V�������<y�¬� ��VH)���g�v5��ѬU2�6�u��o���)�6�����6<�G�)찼*A,��Ўq�WGZ:e��z�2M���eD4/|�Q��t�&�`�8�4#:���Q�������ؘW�,��y���~�J�&�;�z�	����J����(�E���<^��`��\ˁw7��@CA�!��n���}MT<���eym!�W�0�s�
��8=�"��X����}
����tD��[U�a��Xܽ����3ֿ��M�<���.����z�	�\F� �D�(��>��_�sÄ�U�G�bi0y�c^���� �V����~�k����l�qD���O].	��t�Vh��+֦򷫂+y8�^�|@ ȅ;،-�`�n�!$�}�_��9�hZ���.�9	i��*aV��϶��z/Ne�M½���!K��s&o>�W�Q
���^x!So�2+�􀑫F���@y)��x��i #K�|����b9'zȴ�	�..��N-�O�)ԉb�`po�4���[��X|~���x?r�WDgm���r?s��g�,l�"��{�|hB~j&g��@b��)7���=�}��i�Ok�m��!f�|�ÔԈ_0��euB�I��+u��2S�C��i.e�H2Y�g3H�F6S�yp
��r�8�d#rWS�qEpv�
��vD���V%R4�;�z��h���7#�s���#߀��M�:s;��̮�ȣ�%L_�.�V�N���^�~�-b����)\%K�|���ZXМ*��Y�j�K�<�AH._����˂�eč�]��?�Ei���w#�;��okQ�0��a
���=s��މsVI˒ͫ9�	.$ �8����g���M�g���)!FU�BNHr�C�ýץ�z��I���|ͳS�Z�&�XA��+mƯʅ��͔�o<^�� �Ң���6��Oc����a�ս�4�V���k���ɞ(���5 ��Θ[�.�f�<���^IӂY��9H�<`�\�8;�Y���X8���/Mg�ס$�Vn@6$y㎃[�d%z��E*e����k7���ۨ�9R����+R��+��~�B<1����} Ϝ�F*Z�5K3nO��yg�o^!�U
�v����J��.��4�#�qZr[���K�m�i�{W���H�@������T{:��Ǉ
�M �~��O%h�$�X�5����!����|Ml^�/�.�u�nXH�IB��l���@�Gw�!�q�R16�GÐtx�fᄁ}m1*���O�!�p7i���D�����uT�C��Y����̈��м61���a����5�E������I#�C}0{+v��^���f�c��L|�ڴ*C���P�_o�
�AqWlB�ڍ�@M�@�z�ҧ���5R�*���j.��z��AE��lY���_i���Hs3lËd�}��pkڮ�p�M�t�\ Nn&n������Io�+�"��28]VǨOz5 =�����v�nRE���YW����$�xw&��J�׊�ȍ��#ii��de(��zӮ*7~�6Fb�1<�f�$�,ÈuP����yב;[@~�*��:�ђ���n���!����1H�P�qA��K�ZH<R�f�f�t7Ot��#_[��~B�
�����d~�B��(\(b��8��$3
��3Y@�-�Wjm,��~�0�y��,.ӗ�ժ�ֈ.�T��q�(_�����uT��=��4�
L�j S�2�u@�S��bv߭Ӗ~bP$��9�1�ί�_��\>�_��i���&A�d�]QX���������H�e��>�*����Z!�� ��V�����`5���Q�f�^f�@a��>$���Ré�^�!��HY�S�O6�o\��!�T���Y�0(�$ �!����:��dCX�u�A��sH���̱�;1�"����g�3wޕk�&���E=��;"I�2�
�ًL�h4�T�as���bg{�F}7��ƹ��"�=	J��P�8�G���_��i"[�g�7r-t�1Q��n��iN��΀��\P���4] ��x��Z!(��j����y�No����*������#U�a�j� t�q��cK<�Y�:Y�'�Y�_g|��4�9e����
�R�E�K����X�E���IA�`��7SYZ��Z�tn�������O{:�$�j�2�����6hB�'l�[�^̺���k�F,��VSz<AC��͑/�o�i74����� 7�ze�T|wĠ�&�`,���!5CjF���6]T�
 �\��r)�6��xX��ɞr��#ι���7�<Y�H�G	(�}�ơڙh�`N1S^w��z����oYK�@�}��[���Ź�(>����׾U^_�1�늩*w��·���D$b�m�l�����p��t*щ1Ґ���k햟�0a��U�����k�k��3��dH' N��*.�p��dM:�(>�8X��ͯ|�;Y� 3,�ů�	����Q΢�3Ԣ���@-?�X����4c3���agu��ᨱ��z:���F,%Z-��_D/@���f#� �㩔,�����Ԅ��jMe�^$��0�h�k5~����Q�he��Z�fR�(���"."j�t��x�P��r}�'7����7�0w��G�ʺ	� ���Ǣ�<��s ���ߝ�Am�ns-.q=�G>Ϩ��~��Z1�K�%	�o^�L����ԥ�Ĥ_�~�v���F$�$�����_���E�錛¾�\����@�RQ>:~�V����7�N5,��]
����
�KPQЎaj�����y�������l�Èr��� bׇ��o�>��#�8�#�˒xX�E@�dO	���ȟ�fZG�in�������]�ᤄ-XK�9�,:�n�͠��7	QN�i�e��&�@��Qc����'���������3�ɱ�����]��Dl9p���D�&��v�Ҍ�(�v�Iq�����'ViF1y	9�����X!�����X�(����}Ψ{7d��I%ֺko�5�ś��})����=5��q��W�����\�{Yk\��ri�Ě}GM
η�w�b����(����oqG� %>�x*��
 �J���7}#3A�>��`�M��3y4��pQh�_g��b���0�0y�)�r��z�������OT&MD��7�e���Өb�o��b�ľ�ɉ��)����9���7/��2[����
[^t	�AB���v��[ʶ��ڳ3��� ����,�"�R�dw���5��b�����d�*ߣH����g#�_p�dD���8����4��%��v��FD��?p�u]s|9�L�A?����g(��W�̣���+��X[=k�M�xY��A��$�u�k��-m��4RB�$	���(r#ݿ�l�[|Zk��5c�&���N������@ӟ)\��"��lB���9�������&�f̝�qG�е)�~�_L���BJO�~s�!(�e]�<�UOj�il!�2����k���D�D�ɹ,�])n��9��:߹�q���
%��K-A����Y%�(®o�=��Sw��J(�=��ƏP"��&����+��ڜ�L�'}ӎ�(	��$���� �K����U�#_cH�d�w%`eΰ��`('L������� �b��X��*��,v��1�����ɳh��w���� A�����C����.�{�JZ�$1�U�0ZU�C Dx�1y*1�r�
X�b؞[rP�H�tP�ugD�ط}�-.L��絽2�Ҩ�p���V�Hy�x��!z�54���?syh���"T��Η���!j�0\��YהH[_���oS4!�,�J�Z��(M�wap��u�^���;�_��,w'��ƫ
`�����
��t�%�W;�>����)�!���ЊD��N%�e�����;�채���e�SۃFB���uoL�eq��]��]�7"xb��e&O�����{A��eXp>�f냌�Le2+�a��T������xό$�Q���A'��8^C��B�=0*[��B���ײF]Ã׳IF5O�	ť}������(���3M@R;CI��|7/�	؞�nn��s�Դ�r�b��- ߫���qs�������B����p!��g��AAvOb�,V~�xfP�ִb�\�T�Y��wbM�Eo��و�D�����aW���`IѲ���.,k�5���[��\*��쒙��"�"������]&+�	�K�9�zr&ՖP�Ӊד�]	�O�Fa���Z�\��5��y|�����aG	Qɛ���V�0�Rqz��m#�[�@a�sE Q�ML-�}�^��M:�/�Ěج"���j����)W;�Ј�	���[g����g�3F����;`tI�ݚ+'��#���'��ܸ��2�����78��W�$�-���1�ϏNV|� ω@���\	k�.�~Ff{x���jE r��κ"d7"�^,��$�j�%�y����ːv�7���
�b�V�x�^��� 鯩ڙ>���^��`6�����t�)���L��+[�*���.�i������cr���hZv���¤�6|����=�aj��g���v�L"c��?��vۻE5,�����W����~�J1�*j�a%ׁ+̴��-gn�_���0��G�"��;!0@���+I)K�_�ݩɥ���!��G��ˬt�t��E���~���F�Z�qL�f�B#�b�/P�3=�Y�;%�S"�<�>((�'Mt��Ja�
�՘�!
���&��1}�ᯢ�J�C��vyӲ6���^N��"���z��V��Uב�c+���VG����if4w��`�`�d���<%�nKȴ}x/7Kϡ��� 8%�N���wG9��rR?��R�w��Z�}��M
\��y�U6��h'#K滽#�����+=�n�%8n�����O��z��@�_{�eb���	�n�E��:ՙ�-��)C�;u�_�'�BC�ӭ��*�=���Tp5�M�1�;��&�|����m���U+g�؍z#䶄��}��m��rOu�+M�Z��WTY%Y3%�%��b��J�^�g�r5G��J��.0s|ko��p�aqKK&�2����2w�͝|���Dsg>+�{E������h� ���s@�x���F�-��ޢld2����P�i�M� ��9T�j���A9/�LK�[`"������A���
�\Ofz�~�=~,�N Ӓ���F�0O�faBu�"z?T��#YōR��L�71ֽ�Ї���A��4���wl��H��(�:���)�e\��~���>��A�s(1�{I���
�C���.�?�A����CQV�ս�7�h,<�&5b�����r������Iڸ�o��'�m��W�nN��`'o>]�gg�ȏ�2��l_�s(4�z�5����fPĴ���8�aǖnLm�<;7�%㑮�8U��� �AX��|�5�_�����3�9�/�7gpH�@��di ���
 ��oS�L['�^��qs��6� �) ��E������j
���{�=��]9�tx���D�$�ZI���L���f8����kz��6M����M_\�ފl%�~9���زz_O^�X�U6�.9���ƞnsb���[���}û���Y�r7M64x�v��z���͜�,�N�A���X��Mj[����:���T}��o{��>Cf�"Z����O��U�ToǏ=�/�;���5!0/�s�krvߐ��
nx �nA%g�7���$c�[JZ&��}�+uN����/�����8g�G��Ϋ��}�qh�
�W:7�M�m8#i���q����V�.;��줤f-
ib)���yhU&`����
J'�e�6EĚ�}(���j,����*�,H����fD�6�Cșޘh�|N��ͱE	� mκ �	 ������F!�Q�4�4í �<�t(��)��.��h�P\��XO�u�W�(���_��@��$�7|%�րt��V����O�A]�����ꆝ^E��q��W�����N~�_�q����^ABЏ��(�u��%�oW�����-z뛚˓�/����+Iq���6r��?��Y$r���W{OXB�~�2+1>�E�,��F� ��<�5+��"����W<��am�b�D�07	�%b�%��œi�=uX4o,4T�B-1	*�7l��%<{��RK�:�ҭ{'oۂ+Þ� �WB��q?*ؾ~1ߠ-��t֎f�&�h��Ϭ8�V#T�6�]ċ�7+0i9!*�g�Xv���z�����L���d;W���t��R�[�?4��e^� C��r1��ޒf��1./ր��	Z黰n�����։�h �	��{p,������V3|l�l�g��s���gOt�e6R��b�|8�ϣ/�l(Ҵ����;2S�@�z�)O����,�Y�cTb�lw�|N��s�`��tݔl�N9���Ç���Nh��/���t�yg�ńz��]����������B��s�BV��!���tL�=�QSʸ3�� I,��B�fj"td���捘+w] � Dh�O�_�n