��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_l_� (tfvqKT7�߂It����_B��|�/�Q�(Ru؁�Y,F�/���݋ڙ��/�>Pz�	�P9B� ��o��P`|�E����W{�r�(��l���K�x"��� *�-�3
ɠBIx߿ ���K�t��� �vא
���P���1M���g9K�_B�Z��ī>Zvr����ʂ]j���d5&�;�6��� M_aTygR�"�R5�~��8����լ��Ub�hf�� �j5�Ud���h�hX�S��}Ԍ��_�0;��a�9��p&�s�����(��^��Ol�R=7����&Ρ������Q�l@q�*s�rXD�F05D�t'��'��:��+�#`�9I��^P�1����x�R'�÷%��iZ���
���N.��T�ZAo]�U�D8 �����r���@&F�X�طIw.Bt��4F��\O9���r=;�!Ѣ�� 9�%c/p`�h�N~�*�$��Z�	Iq�֧�u��i���aG$�xQo�f�S
�9�!��z%��2���!�F\g�Ħ�n���p�Hf��r:1�f��<8�=�#'�)B��8��%���VFg�9t���<���,�;��2^���*�^HU*�Zg��
�[T*r��>�8�(m�q��#;������-���;RÎ�k� �e]�`���K��2ζ�D���#���D�n������u��0��Ri�����Ny�܋�;�Si�ac�����Zz��<j�kb[�ðv�g�mq	����/�u%�����O�q�����?}����0ܘ�ɫ�!�E4�/��(pڦ:ùg��	����xW���XR7��?�s�3���A�Zͮi�l_qf�cHX|^��ڵ����'��Y���ۊ�����63�OPr+�ȣ�`�?�څ��$�b�%ű� o��+�>��'v�;����b�����0D|�I/��#�#�˚�ԯ/�sT�����!��sFM<�R�:���E���4E����ﹾ%Ŵ*�g�V�ņ� ҤZ���W�姒+6O8�V6�	71�����j��j��W  ���2Up8ErF�hZ�IN.i�I�\�0Ͳ���/4��Ѭb�1�*�K���XJ�?�N�.��aw$˓m�
OSCQ��vm�dP��b�v�*��T'���������Nd��%�v�̸��!�p�_W�ȡJZ��,�	�b�KC)^a'�@S�Oz�X��.���tW���,yV�ʵW՝LE��^l��BW�J���{��?��SΤ�Ѽ�ĦCU���_���'�U�J��m��[�'�a`O�ew�� �q��.�AR�2F9P�%D(�~f��p��V(_k������I�
��M�>+��ײ��+�k�6����K5����_�H"g�� U{xbn�;$�KNϫ���;��\re���.��|�da�q��7�EJ'�&���K��-{.Hǵx�K:`i*�	���ĥ3��9����e���)�0ؓ��Fӕ�u��9br��C�T�j�@���C�[C�HX�����o�� R_s���3Q��]cM=$�M"ذ���@�Z�{��ЄwOm�����ܚm���5�:��R;���|�m����#�Œ�l'�l�t̂�Ʀ�-�����\n,	GN�/���x�F����Ƣ]�߃R���+���ҽ
������=&���r����gY�MrRuk`JN{��5�����3�8|&Fn�_�5�P V�"YҎ3��lB����Q\�i�$�V��Y�R���]`�
u�t����+��z��Ge\�m�k�#��1B�:��9�3᳀�^d��$�i1G�r���Cϛ�7�F�vb�������p8\Nc��*�����N_6�0㶒h`����p3��%A����M��4�Ύ�x�
������O'�-n6�h�I�������=hy�5��=�C��#~���p�m��1V����%�kYNZp�D�]�#�x:���W�-Q�2Ĭ���v�S7-� =�m���صq�z������t?�I�6��;�j�@�&\��˅;Y�
���`nv�4[B!�Vͷ������#��TU��[��W��	�u���?^��9J"&����2���4���g�M�DI��O]�,tm�(�}P��A�1��$��FuqC��ҟ���2n��]/�B�_��O�7��Z>��~�-�z<O��q�a�8G�6������)��
!��@�wVĬ̓�
M[��2:rWW�{iq%��F��0��yR�1�R�&S�>���g�E����]��;����\Q��J�bw�$��M�_0��G4o�oZ��h̬���͠Fm`kBD9�������y��NNɳ �:��+[�-rt�ӘQ��aJ[���=�Gz�$�8-XC� ��)�x a�KVL����O%�E:���͢�M#�Ȑ��ҥ9O���Y>�ꂔ=ƛ���7Q��y NKl���SJP4V��+	��������K�S�ܒ�|�ߞ;��� �[��6���LO��<99���#a&_�E�����Sb*��m����d-J��-�v��8g��'���=+D��X)C�$�&�M��I�g��4����'>����O2� ^����a�p21��s{��q*�G�j�� �U�?�sk�D��:�b���-w3I�T��XE�i�xO"@w2��u�t�TV�v:���	8q'��u�$3sD����I�5�Ac>Bx� \>��C�Ӏz2��4��kgr.٥r��.x_�6��O�x::��Gy��8L:�ܘ��؜+ ��~�A�EDZ*F��՗%>p�~\���i&R\�;���y��kZ��0�?�jJ1���\H�)vsB7�UKe��w�͇?��s$D���ڱ��dvH�S�
%U��S��AFOv'�g?�c�=xI�LkQ�t���,�[��X�^.�e����uب5�b������e n:k���aI��3�����l\ T�`)����9��*Ŏ��L_�jE�yzfV��E���Gb���'+���^!ɠ=SIv���c�����	3�˂B��ݹyp!��"T2_Ȥ�xg�����rnh*����_޸�zH��$c��R5F׼�S�!Jc�� ���+�B�0qZS�2���O喼���Gݙa�� �-'Q�x��H�Xf�������o\ׂA��0�b��"��6$B�1,_������Q�=B�:n��R����!,�A�k�"TM!?M�a��3��C̳����]�5y�V�Vfً�@��X>��H��盔~���Q�%WtH���?� &M�"�{�=`�'�}8gZ�d�p�*T�S.��ʟ��������R�S:M��x��	0��|��`G{���c:�J��=�=?FW����M�;k�0^[�&	T֗4vK7[�p�/'��9��MD:�ύMgn*���)�? ����z��F�#]���&Ԓ=&�{(V�&U </�~�U�*y�H'P�d$�[:{k�?R#~7�r��y>pɈ�|\@�x�������!��/�D
�ó��u6��fz;Xo�G
���#k'�|({�<�w������t2��-�����$>}��P�:����8�v-���53��$��i�|q�s��}�@����P5?���=��V|����aY��z����D��˗fII��#P���ҏ��e�s�k��T�����Wx�G���o����ו�MG>�*�Oܝ\0���q�݈f|t\���e��!���{d�K�*�w�/����Lu ��n�O�,[J�`eO L�`>�pˢ�	�Z�QE�V����;���Fwu�'i���5ơw.Dt-?��u-�� w}����,�Һ@��V�b�V�}��=E�c�usV���I�ue��=���
,o�6�v��Z���K�O�[O�C�k��7����_AA�LF��d�B~�(�&�# ��t�4/&'齆V8v�bD�z�wR,�v����׉ޠ�v-s�'�8�&���1�����}��� b���i�������������2������nR��*�;��F�T����c��cҪ�q���R�Sͮ?�\�N܆a��,}����B��s�b���Z7_�k�p���y�L5�e�px����{���5�Op�c�(���'#��+.[s�c�6!K�)No>�b'�f��u�80�Q���	�fY����s�m��wi��!_�����zo)��Lj��vŚYK�~V�y̢V?������SCJ�u�o���r��~c�4sUΤ;��l��b_K��Z�o	�n,2��F�C���/�h�B��酞�~nWs��t��w�:���y��&�r'*-�q�s���FJ�*�\�,#z�v:�\�^ksN16����'��$b*1+�(4������_��	�}�,ZE�m�E��Wh���F,���_	�C,����.ۜ�4��N�ʥ�^Z��� ',/����*u]�n�
fõ|��E�/��(�>.�-�J���j��� �L�/+��g�H����G[l��N�[�k�	>,�LUh|�E�r���q����!gr��>٨hZ�>��j=Q�9�3"w	��t<�-ra���/�i<���Z5k�����z�٬jv�Z)���� X6G�G}�/6� <��6��0��Ľ.�s���J����(4r-�D�-�n�su��� �xŏ����MM@�L�Tv�9}j ?S�v���XWU��>�=����s˕u8)��U	��jg�\\�-�rCl�%U!Dhն�
�J#e]��W�:���q������%DY�)����4��r�<�8��ʫQb��U���d��m+��Ñw�|3�>��0�����P*V�UdE*
���P���v�(#.�X������a�c�0�9Ibk���M��W#AX��C��������ebZ��=����%9�jC�6�[vPF��&)s{�ƑwW����/�������6�����2��X~�oVX�aD���$ a�+UB������G��-�G��4�f��Y��w����H�/�@��e���F"��xᓃ�R�&/i<�O6�|�	�<��*�M1>ը���Y��nm��_���^��*0��n;��؄f=��i��̱�9&��)��&���H�+^�N���̂�G���A�����Dȣ6�3|v>]^����#���nS
��DmlI��衭đ�g�j�b��ٚ�j@�/���͸��?�C��d;y��BI���[�-?-	{���\�N^P6%f���oɪ��Dϝӣ?�c =��YyZ���]d�!��>��!��HИ}�Rr�JlF�u��Ù})�ۗ�D���v���[��w����F�E���["V�nU2l^���S7;�Y��������H� ���n�$��箃���/�bG�	�Ȃ�dVZy��z���8am��R�����~��,��;�!��S;&d���K92��+s������y�MD{�9u����~��⃐51(/zǗ��}4��Pi��]c�X�v6 4�.��BS��6��28Hܻ�]���бd����,�� n�_|W\lU�J��wr�S���<�l�znL�k��}�\�0�w�r�o��&� ��#�	�o
C�+׉�е ZHp��j��(X�ə�_��/!�J�G��=k3-�M~C
���n�GG�06t��]��P#��	1/�O�CY��2C��g�͛x S>ϣ��(����`=�" �N!,:0��zx긂��O�Y��9C��\�f�Ǖ��l��]HX�����TBủ#�?��p��JL&�U�@���B�@�ч	��"�%:׃����pF3s�ʚ�r!ᦝ���W�9�!��VOM�9�Q;�� ���NT��H+���w$�7(�qQ��*&l�PM+g�-��^���V����"ˀ�|�+H�q��EV��:����!>
#!�H��(;�t��0J)%2�� ��n>�qW7&7��W���t�?fq�Y����!U���HU��Y�BG
�	�*g{0)�;jQPl2����bH  7����$��\���� ���\���K��bəN�;@91'�p�h�{�X���h�P�Gi��^؝RJB�j%�o7�R)�ۨ��������[���iWȐ��ӌX�7�
>�[�"��5d�������qM80��%S�7�E�;~���A��Eb>�$�4=���ٹ�Ag�/.8��F���^c���x�@Ǽ�_d�eUO�]�\�J退[�J�@&�G1��6(�Я3�k��?�}'��{�s�^�(�3��d�8�B�%]�ϕ���o2��*���Q'�Rx�,(HeD��C���b��Za&�ϸ�A:ړbY)aU̶���7�p��$�Y��YR��<;h�q�J�P= �!�jP��w�`$ԷR�ڼ��b��� �q<����ighH���J�}�?:dכ�s:i	��C�<Y��&���(SI�3˩� �6�Ree�fL�soi��/���Б�})�4�W�d�=?'k�NwT��_�e���ҋS`(���\r�K0D�~��O���tC�U���wyr�A��O�F�6s`����a(�Ү6�u$����#L¨X��Vt2�O�A�����nf|F�S�jӔ�X>ōN��4ոj�#p}%GW�ZD5PNo&�-�SB�⧚���\��-�I��S��ZC������j|���3�u�J�����?=뇛y��z~�R	O�9M�<���|��e`����4$aTsH�%�^7��H�S%yԉ��#M�����N#�J�h������U��RJ}���W��l=Eˍ�۸��oDѹM�1�OA�{���f�I�_l�߇P.$dS�D2����]g�.��:NQf�!گ��O��-$�&�L�1;4��sXiL�**��W��Rk	K���7�QuQ	ebw����F�vW0�Y�;j:L��¨�#�U��)���l��H#�Aį�?����t͂ B�=����@lo��3�W��[��1��w�01��*��E�	*S��+DԈ���B�4mv����pL�`��wS���KroI����S��&h�i
��os�P���u��y��bba,u��3�:n���!��j��	,^�I�6	�����:�s����;/�'���N]��7 �Y��l/a�"�ӵ��DX		8v�w�ɿ���w4�&�{�Ds�)~d@��a���McU�K��Z�e�P-/*K��m��-Ji�:��Č�S`yx�Iם5)4��Y%�*H�'Ro\��{������i�G��mA)��q�,K�U:���V�F�����N���Z�(2�