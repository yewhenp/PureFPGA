��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� ��/���Q�?c&*0<�ݸw>V�"WDz�u��AyE����l�4	KU�]zRt�%��51��6�"�g_��Z*х��Vռ�P��I�֯��^�t�d
&�o|0�T��LC�|����[�������И\���|��~�f
�C��F��f�El��џ�0NRKxǃ�����Q\�R�\�5���[�ƣxO8r苃[��"��	�����j�w��y՘�������͐� s������G��}屏@�mM�v�U[�.�����p����|�T��+�D����h�|E�JOAJ�>rU����o3G\�D���Mx�M�]8��IO�ٗ#�}�N�X��Wd%��5�Q:�M�	���婂�z����?��Mr*rv�^ʭ��p��I���0I~��B�\O��q_��dմ�����Id���(����*܂�c0�|+�]����Z��Ae4�~D���T�K����  �'hY1�LB.�};Ǻ�@T�l��i�1�2����Y�S:@t4�x�����XPwK��I֕f^�\�J�$�$��8FT��'�Y2F%f�ީ�?��*�)d�!�s�뼇Y��
"��
r�hJA���W�~_�<Ia���w�c����Wc�N�F*��DaEN1 ;����"����#6��H��=6O� �'��T�m{�}�&Q����*y�Ml�]�%�
T�F�z�l)��"�A�"�(r�T�}0��#ƍ���m��C���:�O@hK�X�ЯuD�T��R�>�E��F_��m�#�%r�;�+iD�^��ٲ>�S�'Pk��@��t�ne_h�iT��� Z�W�u}+�І�j߫ͷ#k��9`!�����&����9k���\p-0A��н��:4�ք)��A�z*�q���s�ue>h�	����s����F�e�3��̻h�@�0�����"�z���6k�ǌ�c?�Z�������� �s��i+�SZ���!�T�w>�.�+(�w�L��`Ih�&��cu���5�p�W���mj���fch����+�)����u	=��Md�+�$m��f��(^J(�(1o!�4t��I>�I�)��@Z��(p��G����j ��(�0�z��U�=C�,aTnl�ϸ���ϴ\���D'c�� ��@Mc^�f�x/eγ������gir/x7�r-a�϶��8�N6