��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� ��i�r�u=
l���bu���mt�6B;	N<K��7�/�f�Q�6���7A� .]�Og�s��K2�)���E�G�:���؍�2��
�?pO�x ��2�-����No�����ۉ�j��QP*��e��`��U;��F$�o�J>�^���X�����x�Dmm��ì�\�ٌ[J:��CRF��8�r�ܡ�=�z0���,�N{���������Ȉ�!�~R�H����'���]�0��K���-������q��R�/��+�m�%��#�<��0(����F:��ǵ�c�JU��*�(,)�`7$A�Gd�"3�8P�杸+*��RUsF��A�C���<_��H%[ɠ��4
�������Wp���7��][��-�E���a7���W+1�`	K�"���&y�B�����`6H�˔�.���j|�o�w{��'���p�(���:"(���%��>�'�uR`ߙ͖��ΛK����o'p6pH�^���A�aKFRT1z��v�\�>jdq�H]�c\�ŽM(.x���Nq������$z���9�P�w���dB��p�q���5K�+��_ �i>ǘ_M���\}�Z���+~�E�?�F2��|���"[#�ӆLǃ@�v����2�J��jh+����ޔ�Eq�O����t�GA�iT]b@��Y����ip_��A��r�v�vv�	�#��Fό��@kx;8.+��xHJ㜉x'
�.J67C�)�����,�ft �O�NQd�w��6��R�ק��9��ހ�y bL�s�M
\-���� �}d_[[���y
���̒S=�ɯ�qȟ��0Ȯ\䏤QR<9m"	�=�g�u�-��c�_<dk�����;V�V-S�îTc+-�}��3S_e_ED��nђ�һpY�{��:��i�D�([&�=�B�ت0���{q���2�n�N X��!P�5t�^EH��t̸x�	(�L���4��᧟Qx�.;�ߊ@&���3_��LOz0sn�Ł����ݤ5&�w�t��P�W������G�G�M�(��H�da�=�tKVr�p3���\hL2n�3�hVE�/+E��U ������}P=.*�/�d�x{�*���Z����Ivo��|�Q跾��0'���f^���a��.n���PU֘�|*� jO@����|a9,����;�H��?Y6ܘh��{q�o�D��鷝��T�DU�$}���Ĺ�����w#m���{��Td�����VO�{
\f:�a��})0�J��}��͟ }�d;�N��ξ�Ǚe�h�;�̗9Q��#2d4Z9��V!�i[�Z0�jP[��11�D!*��lB3�U�JQ�)��_��~4��NF�#��%��"	ƶ��L|I$)�!y�l�\vR��uݫoGnm�\p%Z�b6l��¬*�nxx�I=~�R{?.�w�Q@I�-�6;� �7��uJ]�c�O;�^�K���+=�?�����d-�M������0e![
֣^Kw�qS���GJ�;h�H	��l,=��=�Z8V��j>��4��
�y��Y����c���>FGs���^�.}�B��r�~L�IM�����S�������<��1��-P� !U����k4seQU!ٞ#܀o�};����k	���ce5����o��o��X�ϯ�
�Wټ�3�7V�tI���k�j�ߟY�׊�$#zǃ:4n���W����'��q���l}B�W�@��ǖNV����:��-B�`���A�?J�`�D����$k ���W9y�*��j�E{)W���9~V��n��fY�WZ�`������Ly��f.P^޾�m:��)�Cym
�l$Q�P�i��HJ�/�g�q�Lh����&�4�yBJ��#��^�Z={-�Xv�}��L+��+���vt�^[�C�b�c��:e2�
32E;:�T�3-MD���yqE�Z���o��|
�m	@�`���Q�b
�����8�;4���%���9��)$j�|7bd����_wt����Aj�����ě�cs�"o��f���w���7�`���i�V�l�8�J|��:�{`��k�7�ES���4:���Nl��BÌl ]��:�^-ss����k�����!I������u��7����y��Og�-�HA���a�