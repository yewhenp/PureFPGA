��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ`T�}�w7�ɴ��劂�[���U*i�:����T#j{2+�t���.�h����q�ˠ�h��ͻ:��#&�E�њ��6S��$�}�fa���r&.l����M�^KL��W6��<��:EЄ��1�܍�����
Ѹ��> �DKɦ�Z����yU)�(�:p�Vx�m�C>G��l���>��(ւ���_�%D3M���Վ仐�wngRR��Fo&}|&O��<M�:�k�f_� ��SE�K#q�><����5W�����X��D��^�VW���Q5Y}�{V5����ٲh՟�¼�����1)�b���(]����'�"�唼|�#���Kz��9�RL$��{?G�=�S���݀�m<(�Ijl���ʽ�$%���k��
�f�<��^0��#�`�� �9�H�s
@.�7�0ZLe�o��Z����.����Cl�zf�byŪ���󬞪g�#$�H���0'��8�e!6��֊�����%cdu
�������ϗx' %μHJn�bݸ
>�?h���69�H��=��o�x�vw#�H.1�|S��ɮ!�^����j�V�š��
�Uw/>��uc%
0�FY��F���"\ԟ��>b8���S��ք:��K�1��|�'�j=Ϫ�t��w�Ke�&z�!)��d�O>��I�]`�fqW�;�����v!��i�R?���De5x r�xI� Z�L���"�<lx/>[H�c�,�S��D3~UZ�I���у=h�m?�*�H�4��-��Ԛb,d-�$��9��?�C^^#�0�OP�.*�u<�cRWO;M�=f:����/��i3��3V�T�,�t7��s����m�t2@�s��0 �a�gA��d�m��� �
Ig��&��bXR��z��B�gT�{��IM����C���mPϱe��C��.+y'�0Oo�4�����Cˋ)脒wY����w{�>ʞ7���*c|w�N�j-S��n��K�Gd����� ql��o���SeաV�9Ġ5mD&uGd4M�&��G��3����I�ꮦ#��a`p%���I�����^�v���P0r��K�^%c>����<m�&�Y~v�T�Lܗ�N3�l�dI��6���-��&�����(�SD"T1��etE�<B� ��̎ۿmE!F��.�s�_�ubb��\Fk}��4-��U���SU�n�{́�;Ay��p忈K������g?݊%��m�ηc��]���,\��3s�g�b= �ح��(�~�Tw[X N�jj�IJh�*>���	������WUp�Lh�
�}es�Y����Ug��o�*��k����E����F GXq�AkX��..�20];�h�:�oRva:�e�����[qH��B��k�R:�hhZ�:�(D��C!"Wild�vxʏr.noer����D"��R1��&E��+�u�^�*����a��N߳�_i��}��[	z�vL�7-ӷ����}�1󃩾x�:�8�~c���#,�3/��S?��dp4W����t�Q�M��;�)�M2�j�a����0�=�T��tn	��.���=�K����o)^�#�r�O���G�jg{�s>�VK��B��[����>����!���,״�&���cܸ��l�,(�H�����D%LE�p��,�}@c���<Iz��!5gx�<���N`���nYXmq��2�EI�9�Q�:XωdMY�8�ˀ�	���@&��$F+k�!u�}�ῃ��ݴ������T�}!k*������;R������$��^� g�6f�=��ac���d�l]ߤF	�D��(!8�5�JZ��cEm�ӌqtU٪)o~�!��IF���1s�@��θ�%Ū(��֋��k�-��]W�W�&��LϮ������ UN?c�MIJ/��X�[v.�ZF��Bє"S�#�Ug���а�j�{y&�;�z�<YA�{���G �Ƕ��ؕF�/�!��j��e�(�1�[�%+!���d�;`�V����9&�H.$(�<�CE�1�r�?�0��ݦ���К�P��(Ff�w��<�Q�s�e*��-�7��Ot�C���I����rq2��?C�\��K�1��d����e;	��.P�T���B�z�X��P2(�z��2��f�ok��f��x�ei��K��}NK�J�oQ�I���Vv��(4��;�)��V~��D�YRע�2�hQ��Ue�,!M����
�������a	��2d|�)Ex�
��s��v�͆ �$�~�ۀ]L���Ow�mv��9�\B~"�6���%׋/���yS���LK� ��0���$�c����A��@�LӇ��H���t�詝���s�c���ODz����~ �%SB�M�G�+z�+d���(Fs�2�%<*�I�}��v�� TIO�P9�-��/@�/�,��pr�JG#�cm4gEbp�����SNT��]�Ǘ��]�
���p�L���ׂ;��9:.�i���-	���xv=\ �^fmS��3k�#y�!�m��E�D� z���z"�X�3��Y�w�s���=~�L�y�z�^p�:���S ,a3 ����b"&Bv<-/~�%�,"ɄJ�;����jp�b��?CF���`�� NJ�	hy#"J&	��EА�<�h�q�
�p�L�^���O��nN�U݌���Fe������
��@������M�G����4��^��;�h,�aI$dҺb.A������˦���/��u�Xj����(kt�l�?Q��-�����	G/� .-|
���l�����$�C�PӍ��BW&�%��7�3�$ēy�2�蛛(x�ʛ�I�9�����_p�uyǮq�#�D?8��2����I܅Ԏ�UE��	Li��_��Jމ�Ü(�H
��m9G�]	V�I���1�a�׶D�!�|�;�	B���S���JJ#���s֣� �;��2�Li��ȓ���9f3�ؘS�N��0k�-��ڙqJ��λ\�-�^G�*�t�S@�"���(���Q���n��.��ӛ����'*�u*��h0�����V~̃}m�N?t/�������u��:�ӂhD$���6���.���l�7S��Nhb�M���x����X堟�?���c��Y�~�	�N�1<�(�PN���k�mK�N~�p7r��R)%��%��=�$}��o�*�"�tNAz	gE��Jq�P�V�T63e�쒮H4��x���O+�7�8���Sd��������,5��^޻�9�
}zb��/����_����+�'mCo���;���[�e���\.��?�H���9�\������?[��+��c4+8`��(`!d�ɞX�:5���������za�����XL��[��R�#�����x>�Ǔ���� %-7$=m�q7��U�3�����Wq%��D�v������O�$|x��>��������
ց�̙���xz���֛/h�]�h�G�v4�$U_0��Sd�c��hC;��v;���s�g��_$��#
k���\9e��.�Q�zrC 8��ʪa��/+S�!�+���݈�~!�&�%<�7s�|�#�k�UM������PH��=u�(׌O�v�� �ㄌ���� �˼���<�bW�6���i�&�5����|4-b�;��Z�	�)r��|�5�Ի���oa�5X�lg���S��O.Y�ݴF^�|��B1U 5�xtհJ�ئ'�-�;���,�9��#�N�o_�DM)�7j�37����Og���%�/��G#{��Do[�8��Q_W���d�m)�ggEy�SbL� pD��Q���8辂z��U����N�P(���v�H��jҟď�j|P��ȵ��h�y��~ڬ̣W�S��{�S�JG�i��Na�y�Vcna͏�q�2q�dZ[Ľ�?LgeeM�q;��}�s�F�stEK�ER-M�G��{���^�A��o!!>O���C������ř�� �na�Q|h���E�W3�4X�o�1韢����l{���/7�fI�JN�B?�'v�=d�yH	bpB5�d�<vfz��͵J/!uh�G9����)N���.�����̫WE�������8�w�6�r�g������D#a�c�om�鍝����}NT}/Y�b7� ���i��a]xP�'.��F#�Ԡ��'U��j�<6�M��;B�b&�1�I���F�3��\�WV0��C��Y�ҹ��$��2��rq��w]���$z2�_0�pz1����dC7 ŷ�`���!��<�d��]�h [�����Ģ�$���Ȣ��E��Nxu�Qx�d��)`D�� ���}�f#�0���&��������Е	���ʒ��ٖ��Y�!���P'��"s8T2	w$�L���u��0>���}�(&Ph�&�Eu���ԁV���dt����T*?�S�Z^���*�8e ��2�������uj^ey��Z�F��д���Ԍ}�J����vh�z�똡��z�?:ӑ�a���L�,�	AL�De{�bdSI@�^��(�s��6 �"=�l��ڊJ� ��"ԫ��� �kh� ��A�ޭlJ�'K�=0Q	�=����n��7>��.(�3yV)	�O{�q}xy���ծ�Þͪ%���@����os+�'��3�_{2��x5�W�v�BfJS��KD�
zq`�]��ۧ�xk`$X���z�S�^�A��h߶����0?b8r����T(]|��V}L�{�ݒφ�u�Y%�G�*��I�D��P?����6K
{���P}��)KX2Uܰ��g�dR�?����"Zd��*��WXF�V��̀���,�
ݩ�:�?M��8d�}�S�ܳ4���z�ql����+�D�[Y��R��Jj̅������8��d8[Q�w��ُ�x���%�n��?�Ղ
�7d�h�u;05#U�h�P�]N����՗��Oh���_.[�\�5Bk�>�]��e��qU�H��kga�3o���%������B�z�	�z�y�Ú���6��lߚ��*Z�}��rW�/`e,�}Uw[�Q�����`��`�����[�`w��t�5��LyPC��j!�E�D~��V�S@����T���S5|Xc���R��+�F�����T\�.C�VH���`TUɀ�|�҄Ec(&���]�"�'u�k=+��������������}i$�P�LB����&�4ְ���Q$H[���D�40#괽'���U*�2�T'<�Dh9$���D�`��4W&�8��Uk�e�V�p���δJvw�L9����]*m=H��C���_�鲑Ҿ.f[���[�v�?z�	ˢ�H�rKx��:2 {7V��*�ap�b��-�,���Z���!�W
5Gr]Z4=�ڕ,�V�OE�Q��CuQ��T���M8Kt�1�WHuvh;;Q�� +��M�<V4�����e�G��lUX�v�?s�Z
��!=�*�Ϙ�i8�+<���KI�7vD�R|��(1
N���L��hR)r�\b��ky*5�r��$��^\I��o���V��R��b�O���jD��l��o�S���L�k�%����p��A�Zq�&�O�i|�E -���F�,gS��(Չ[�����oR=����n��h�U��8O%^�Jdq�E<�bh�}Pb�ڕ� ���0�,��8g�l�\��˶�%g9s|����)�m�C�+�Ec%?�HZJ���ͭw~e��l#us���jϬ�'�����ót�@�Yb�Fg �X�F��K�	�� t-�^�V{"��GG�B���)#Z&މO��$}���*Y�|�+YN��O���b+��|�X�E�j����շ�'R����O��7^�1)'� q���M��ӝ��v��B����-r�j�5�O���V�,�bY] D��0�eБ/�_�r�U��$�� VT���Un��������bZ&���Y�`f��<�/�L�����ȁ���G@ï\���`��t���Ϲ	_P^��Q�eܘ�f����b*5�qI(.H�n�a�;�+|m�u�DX�8�"�t�
�X���ؙ!�f�~���e�W�Ur��R����WP,f�n����t� ���P9Ud+F����y9T����GOh`�����I�
7�=�_F���l�f�jx-����^���bw��������[�sX�ˤ!�2Q�īӅ������]B�D��z�dh�"�Q����>�2�#���c�ah^�W�� ��!G��ݣs�u��P���i��2���mI:˱����.[=� �Ыa}4K�"d���;[�9���P�R�l��@�Mf��w��G��Y�0���E�ۜv�d"p���&����8�J�)	O�%{�q��?�������b�|Q����ux����Y�Yc�GAЍb��-��|��<�(܄�,�{�z�2��>q��i���	P2蛒��d�~^���+e'�Wb���Ϳ.��S��9)�6J���`]�3�S)j	��[�$7�s�X3C��w.�'a^�q'�1��eW�9�����ؼ#�u6��}�Ƀ�xE�\z­�@�'b��BJ��#'Tn�V������abf�"[�/�t �뢃p��y�)O���kU�hD�t;2�3��BVbSX"����8G)�
C��RO��?KȬr ��0��þ ��Y����yNc]L$�#4�����B1F�E4ȇ].�>R��	xBLgi��R����� ���w�6���/�N ѵ�Lm9��������V����������޴X��+$��9��ޢ4�X?�->�7�ײ�&x�S �����_Xp���9C�ȼ�% ����:H;�`��MB�~�R��p�����B�,8�HG�!������y#ӴY�{��?1Uݍ귾^Al�{�����X�{���쌙�ɷ9��ţτ�E�0d�	�p��>�F��, m��E�����ǉa���M�Pu�������VRht9�]��7��<�
���p���Wx����Ig6�۴T�#��Ýl᳇�Qo;�
I�A��i^���H|8���.�3��Gd��rJ�y$�H*��o��!B	\ܥ)��\��N_�{�{r�&�@F�1��� �S�JƮ �&��]u�<� %;aW��)ϫ-~�p/�'u�kNf��^��!ҭ,��RP��aj���&�H����­HQA:r$�a�쐆+��|�������l��p��h�d'}.7��n���߼�>��@�Ԕ��=��D���YL� 56U����8d� "HєRH-M�i���~ˑi����]�{׊��6����Od0��0^΄|rM�rm�3W�wV��J��d	D$ձ������&���E�s�|Q!�n�;��w�&L�p�qԿb�˹��zo�� |5�$���[�/���7�� osX��ڊz� ,����M��s�N����++O�S ����rH^<���\<hS0�	!�w7�	���X8�&ls��@�"���י�×q�^��E�STn��pv�cb�� �����UXgu$�:���Mֱ͆T��#?����)�y��+�,�(`<��j�P7�\�N�T*	���`�y��&<�O����*|�.(
�]k��x0�C���y���0-ӂLt,���r�TDn��ϛ���F��&����fJF�2��T����Y�0v.���y�uȨ8�HT�V6����_RZ%�X-�/\m��	2�̰�]K�����Kiv�F[~��P�IW����.��*��I]��`m�JV[���9�M	g�۴�fљ�����-=����3�4�ۻL��	�n�i��g�y#K0���h�D�VCs���2r�_��p�i8}X��~b����qS�'ޮ t\�S�s&�n�����v��9Blf��*򉹆�����_z)�+^�{J_��@<���L�vX�J�D顎7�aƵ�3�~��A��=�Fz��l��?�#p4����#_�.����:2��o�@3����G��,N��N`�10�jH�����2!��Zs�Y���j�N��oS����埋Y6�ᬝ��tɳ�����b�� "�ݵ�\�9]��v0����0���9����/��x�R�3��c��q������K(�yb�@5*N�O��E�s�Z��rRD�nl��]�I�},�^K�"�huդ&ys�c��E���;Wx��Lb/�yޮ�6Ҋ
���ո$�'1�X�&�^~�6h�$����2�r{��Y.��DL�և����g��%E�q~�����ͤd>�mM�^��/A�7��� 8�g�ĶF���O�s���7������c+��Q!�S�)p]�.���]�F�81y� �R�Sñ�ר�14嬕�z�u.f�w}���M3$5�Jw��g�­ɾ�S���qa�n\W�0n���_^ɢR�zbK���ɥ���Y���Pߚ\��E��|�q��Ҋ�t]��h|^���~��_����� �� "�
�
8@��Є�h���!?s�[ʧ�,C�D�̟��3��Cq[�d�j��
��G�p83��H˝�d￷�Bu�94X����D����q�:@'�A﫚>��/��9��J$!�+8��9:��v��?s_�t|K���>y2�����s��2�!7w9g�v�FǗ�u�m$0*��r<��Gޔ�1��uj4�W��6Z7l?s[?)�Y8��9�HA_��5Vq��0K����+2��
^�n�c��v��ݺ�2�����!'�����bp&9�+=4�'>׵.�f{-�d��W_�F��qخ���C��$�\�_�x
V�
2b�<K��h��ʞ*ز��C�(�;�u_H�*�qw���[s��E��l�G#��q�wS���@�~r~�	��n�5
V��fT���g��$���[���śk����?���'���R�D�U
��!�D�\�P_��(li�I�����GG@�FL]�|e��0$���Nc�X���l_������W����8����϶yQ+1I�ԐE�X�:�A+z�i-*�R3��b�|t���S�:�*Q�d��������_TpX�H��v��ξ�[x��,f</Ng,;kе|`�)��OL�J�0�V�jyVc�|��h�5<��~ v�r��y����T��r0�JJ�n������n�k`m������Y�>����"���\�h�s��YX���׭W��u��&���0FCR+���^D���к�b�^��?���O%�}�_�#��p>����� 	OI�Ӟ��~,Q62���vbéѽ�ے���B�,����6�+?�)�v����Clq$�}�����D��T��9�4�%ĜR�op-���k+��C�u��G��:�y
�3�ɦ��R�㤻8�D^�쌴����/�ǁ�$~H��%����D'~��A���E8{��������ѓm�X�*t�������R���ؿE`&����|��~��=;�b�%��c�"<�;��-W�۔U��duC`ZL^L�E��c��0���He�0 ���n%SR1��@V+m3��Pi4{դ.�I�p�ɬC<he�xAw��C��#��_��yq�bn�!��sF�hلӓbÛJ̬ �<^o\]*�.)	f��w�H����Ǐ�C����.w��*�|��s��"M��ut��M�{�Tt(�䃒n��D ��ι���m���*�ک�:� �z%�`p��g+OXF��5�a�T��1�����ջ�O��:?�E��Nr�P9�N=:�� qK`H<�P�	O��Y�~�����(�x��}YA�!-�ܑ�a�n�B�t,�W���E*7�s���Kd����ă���<���_Y*c�'ykI�vq��2��c���g�^4��^�J.��%�5V<|��pQ�	H���;J{��k�@#�j�22��$���@P5 a��U�Zs��Kp��h�
d��i���G�〯FO��93�ᇐq��x�D���o�b�����K'�fa�ס�C�h��h|�:���`�C�`���5�lgH�Ad�~�D��8g�a�-��1ZL�v� xI��t:��҄�₮�]�dR��`��ڻ�k�k)|���/��w�����B�y����]����.|mԑN�d�	���{]�gy����H�"�{ Tt��E�6:��P��/4��PdN�T0��vo�y��w6�&�K���F&,L��������)?-k^l��[�����6Q�2��zJ�������*��6��'��z�OǦ%��R�C�ys��T�Ĝ�C��J�p���GqX�0��j"d��J�WC���&BI�G��W5���FwG?�C�9�(+��E����	i�_���RP̚~v�վ�C�� /Xq�\=C~8BbS��Ql&��^��ԕs��(��f�7�څJ����XӎJ�6K���@���'��N=�_�L��#;�#�����e&V�۪@�ǃd]6��i�Z�t�e^�?��{�0�DgRrj-��x	�*30�K�"�t�w�*������;��� ��o���U�b<
T�Cp� �c�	��9����a�pC�v�n��i����8g0��zOB#z����Ҟ��k�"��A�&f��Nצ����w��Y�/��1����9��'��d��&�NZ���/m`�����Ws�(w��҅kN5>Dy"'/�X+2.mۅyH�������)
?���m����k��;G��	;��q����.��q�WY�wu0y������K@׀� -��/�h|�z��m=`� ��`-�[b�]�̈́]d�����sI�������F�p��_~٠��4��q7> \�w�H_Y:����!�>/����`.Ŭ1쐱����P�&;�+��ӝ�0��~a~^V��v�ɝ�;�t����q��U���[�Xdx� �?vB�O=��ë8�[���p�+��?F�0�i�F ~+	�輓�XG�̭��]�� 	#�+
���:�#^�b���
�z,��u�`O%���c�*��*$JRͧs,l��a��_k�;M���,�����Hw�ʟ�yc�}����Z �J�P�CSb�y���3��s��%z������7�Q����3k��q�`aB�(??�7������[��˾Ѡ Y�� `H����P��Q�Yc�^������(����U����C"��J�kh���O�Ah�{���/���~���)���fR(���i�G���s��l�o�>$��F�|'�S��/��@�j��A�Ja�tx���� MOHfK��.�\\#.������j?/��k�LZ�LW���@�QLum�{����C�w&���?k��ȭ��HD��0+�D�*�N<H��\4�Sۅ��S`����)��P@�X��vE!��6�d�_�{�����+���2�'$2!P59���� /��}�{�C6���� L���3�CouHUQ�D@��n��$#L"�'?�Ζ��V�����QlMBOmRQ������0��j,�O	�x�7+L�ˆV~�V�z�Qa�PSR�V�.� �mOE9bV`}�f�S(�W������� ��+D������vE��0�5&��uj�8�E�/�A|݇,-���ԫJ>�^�~ng�w��}�Q`5w�����	��\OO�q{�%@kE6���cwu5�]͒v��*�U�X�w23�7h%�{�1\���f����|% �w�^�09M�տ��q̻��Y0kyF!2�Mk����P��w�*ۻr�R��-�	��`#p>�7Y;6�ܵ�97VtI�7Q��=%��gh�����3���g�ֽ���u�GU�M���(��$:�\����q���E�b��v��F�{�'C�����s��N�����S�~փ�������Rn�|��
^�j���4Ia+�R�떒�4�!���W�xٺbɶ���*�6�-v]��Ja�
/�I���Պ��If5�b������"��|EԷXZ>N9Ϫ����Y��4����򁥜�N�P�oEP�4��zXT�>A�?I������k
5�H^�����3߽e
fZ����{��/�j��ma����'Ю%|��]S��4��9���]�W���睘+�|�G���~b���{=*��u�Ɉy9��ll���PF�>a�<U�D�"E}YC�w�����neu�=�
1���hMQ��3%Q�K��UK�V�xؓ>o���%��%ľ:v{6�^���������|_u��	��k�@��6�'�g�/':��p��/6s��T�	���!�P:����[;N�V~IYuvƮ�����3s���<����RTWQ`�AnV)�6�S��N+�V�W���M���v��SH��*9k�X�� )h]��2��6Z����Ajky�)�,�e��P��G��Y�����4WF2,GQOF������@Q��S*D��A ���|O(���m�}m������E���3�&Ӭ��r�tkΝP�A�%4m��̽�j����Ǟ�
�9����Ri�bI�=�f!W��G�+X�1��o��<	�̧Ә_��|�$�zI]�:~��N�e?Xߨ�ڳi2�i��HQ'�Ox+)d��V5�ߑ-V�[��d��FѦL��UC6|;��ճo�ʗ�A��e=�w L
�����G�H4�ue`pY� lB��<ŵ@�a|�1��F2dl��91K��q�'��s4U!�%��d��[~D����,}3�E^��N�
^wӡ6>Nq�� �&-�KQ}����'��W2V�W�sD��Ν�]��,��_�\��I�K������^?��q�j�R0)7}o�����{	�<�;���+S��惋X���'�ƈ�{��Y!>�50���d؅�饐�^>&�ǘǲ�)�`Ɛ`��ѲT4�P��V��;�,�w��I>�%er�-ft�u����+�ғn�	MѨU�uo8��ʘ���-:¥jn�������5�?Yv�ZG��q}��n�-o7�r�L�aI����{�;Y���	y����|ƚ��8��v�[,��Ea����4��Y6}���cz��~�^���R�ױ��ۜ.�-vK��t�6�ߪ��7~��_}��a�����W����d)����~��>;��,A���K�-�8g>T)��N�B�YV�ѐ�+O{�b!ϛ�O��b��606��tWp,���8P��	M���0fp�s�J�V�g�yx)�voi���6�_�!�Q�A�I�3����K,��S2�[���2���l��~8���3� l�#SF0�����7#�e���?���ACm*�j�I������02B�e!�jټ׋djm�� �P�����ǈ\�]���5�iTt@�xJ���*�9�%/�*栋�5s�}�²�D��ѫ'����8	w㙚"T��=�(�j�o�"(Eص��-�J� �@��j҄G�K�E9�ڱ�(i��|*6p7���-����L 6������?��_���^m�����y��~����/��KUg�2�Z���\4Mf��r#�3��Wl15��g9�Z ��GD�T����_��+<n����,��tB�g}?�B��7AR�x_��(a��u���w�Ra¨�|@(�����Rȁ��jQ���{Dq���fƖ���d�V�VT+%��k3	K�N��p���!�C-��=�9��6�w���RY�������BJj-�7��d�u�(|�&�P�����Z{c����ǂۦV/���x�;�����9#D�/�T#K��r2�Ut(.0�9�!�5!�� �S��FA\�fzN��M��Iu�xfF����������}�@�����a��-�~:��#�W9h�m�#�E�����1/z�9񒥲��"��f�W�܃zP� 9�2@Ͼe$�GO�ccӿdN�H��Bg��l��0�L ��=#J����^�P� 	KKq�ܝߣ��0����P�E"r����|`&���O ��5�����FV\��-��%y�IB��ׇ���⇴�2%x�2h���;_�a�r�g�������r�)��g����˫" J�@��m�n2HܓXRa�ۋ0>�.��ͨ3G#À�8������:�a�1!ٰu|I0��!.Kߥ'�+���?I�SMH׸;�	���8=�<���
�S?���~���Mn�����̾�Y���m��\Gm*��"/|O�U��x�-aA����f�!P��06�� ��h�.|����3�ڝ<!De�o�Zh�@:?4�]�6`n��2��`,A7d�Kt��L�<²=��\d���䟽��F�f뤋�]6��U�'
�
&���)�-��9���l�Fy4=�Għ��c���1s�Ғ*���s̛���f����h�N,u*�M�O���8�S�{{g*:)K����9�]���B�ȍi؊#@���ĝ�)�e��̫�'��%��1%u�ֿק�%%�T�`MEfP�/�*9�Q� }~I͎0����b���<��O��b�"�o�/F�/]������¾X7��j����]g��j<T�A*�w��;�$,��U}͑"�(! �*c7��p����sj�"uH��цR#�ooף:+���So�m�Σ�k��|?	t�O��]�"��3>=���b�Z�h�ϕae=f��&�v�����"e:�5��?4AB�(��-U  ��Z�nv@����oh`R��r�;�I�!�_r�=f�$V�>՟Bj���Q\0��G�!5:�G4{79[��s'f(R�]�̔Rt�w�r���W�����
�+P6x%�e�G,�a�X�"�N#�s�`��?�f[�� �IE�n��<�/4i��l�Dw<��j@^��jT�Gd�����p �7����Y��)��APR7:��M./&%W�pX�N�����2uښ,�%vi�LG�_��>b�	)0�TM�"��E��_�= {t��d,$"2�Ow-c((\����|s��/I���8���?*vf��ט�ن{�8�z���:��0rH�����;m�Ƒ��i�{���RA,cv^��ǍF�+�7��:<NL�QU�����Uq�s��
Iq��'�F�1��[t�I���1
�6oٙ7X�v�q�6��LZ�th�m!~�\Zl�)���GlH�%vǬ��k�õ.Q�a�Q�{��dݗW<\HR��&}����1K�m��lU@=@�s.���|v!=�Q��J����K�|����;,\�����rA��*���n}2����c$x�[�X���K|���&n+�*_��-�O�>�x��S�U�$���_���y��e#�:���z ?)��8�mQ@.�v:���\�����g��r*���]�Z�+#ks·G"�����x���T�C�\S�3_f�#7���ľ��ޛ����a@���%����'�L�zlqm���Y`c����yjG��S�Mc]��9�b��p�Ȋ�JS�f���� >y C;��ob�B\Lڟ���#~		�B�]Y����[s���B�G�^5�a*=ŚG쐭��Ao��#%Y�ü0x�)K�&YL�
�vB|c,��/�N��ƦVr��`"��_F�$Ŀ�~�1���
�T��P�*wfD�:�c���\9H�_޺�������(�������W%J����4��O�D�>�Yf�ĥR�L]Vځ,j#�ή
�v�!^z���<������JV���h����]�����=�6zy��b�\�b�������7�S�?3�	.6�;�t���m6��s,�nB�ޢ:���;3`ὦ�7��bO�-YẂ��8 �c4x�]�a@/�y��Tp�t����0M|���	}��b�(Y>\S�o�����h�h6[�Zvc |^���採�!|H�4lŦ� �>��Xv�	rG jE��йVd��')��N��ܗ�G�j�F�6B!��䖛���Y�ҩ��ǱѯdO�t�؊W4:�h�V�	е�?*e�ޞq�%FhM��'�u�O�ܱq�R����Q��u�8���������Ϲ����g\lhjh�1
�y2%2�^����=��@XŦ� ����z�}Hfu� @�D��,��֖sU�`<Q���o�O�擬N��ɸFf� 6��S�%G���pՅ�*.x9��2F��-�ɰ�����PdS+X�}��_��,eŻ�V,�X́�d<jė����+�& &�SR�w@�ҹm�P?����{(�&<#qqn��s��g���bl��Z�Ԋ�c2�s�E_s}!>�	B�w8������,�
��VA|'l�?��%�7a���qe���bs�X��$	�f�Է���Q_RPh�{�9�y��?Fܹ���L_��(�����CҺC�p�q�<�2%�~��]r�$�/_��6���F�HB�P���\G3ϖ0QU�)�Еצ� �E��B���F���ϢZ�r��ȫ<g߿��m:�@!��7�:<O	ˉ��O��qW�,è���@�6f�,�ۨ��u�c2�h���I�4i�%���=A�k�b�-iE��"G�Bޫ���;��4�	��p:w8�Nh��	 ��	2ߤ�Y'�zc
�L�/yv1�����#7�}��LLƀF�v��%�,H8 ���wɣ��s����60�P��j�#������f1i�?q����Z:D�+8S��.*m�^���<���o�|�}�i,�%ޖU/��p�~���B�' ��܁����$��� �>M`Ek�ե��y�	��*R7:�)��ڐ������7d��6\̤G*���F�}�}���+�}���3�Y����z����u
��[�Iig�Z�<���t�b.�+�ĵC.!�6ơv9��ESx��Bd�S��(�L9(	.�|�f����I�x�se&o��)&_�;����zW�T	'����	�M�gWҒ*.���F>����A�X/��{u����:��@VM�KO�mה^a:�6_�.l<W��o��r�I-R?+�m��ͥC 3H��۬�p��m��s��H�(o�������I��6l&4�(?�	k��Z3�������5�+�U�u
���΢�V����JQ;���X�)�qw�-��;㨩�� !��J�M����ڐ�>��M|T�`�U���ps>����2.b����s��Ā/Do
YY�e��	_���k��E�BC�:ΊU�Q�tT��F���R7Q��/p����ޖ�>�!�[X`ۼy,��T�q��Kb�C��|9`@�+�_�`����W��j�|�$ ��80��HӬm{�W >���Q.s�j���d(�39��ڪP}��_�mk���N�ZZ��_=�s�t�%�����q�N����g�ඏ �P�vT۠�.�>���3�'�K@Ͼ��:��n��`���	s`|2mGUc��I��'�}�c�%A�T�(��1�4�G5�*��G�kF�}ܘr'7���BF��28J���h�p�h��ǜ��w����B���h��u.�����Tۮ���iy���t~G�p9�.hY�[�"�uc_�#��ǚ�6Ǧ����.jV�k������Ŏ(������6����p�c�B�h��gs�F�kY0%�X-�éY�ѳ��W���N�M1CC���#_�gq�Ct�=�n�/��������h�m��V��}BZʧ�M�h��]�4>p�xO��G\6�Z��:-��n7�X��E�Cӎ������P9�IL��_9>p>�@u����ZB#1��r�sIƪ��dm�8H�k�	=�.�.y'�S���X�L/����a�&0ˏ�����9H�}����v�s�� �gn���I\ S?#B1�<t�94`�`5����Ձ���}n���=����4����:��\#}��}��y^���T�YR�ً�O8��B$���W�)Q��:Oײ�LQ�D٩%H������<��$�3�ݜ�}�>�-��ϬRÐCe1c� < "/����h�-�|J3=yV~��
�;��:ß=큹-��[�r�Gm�%Q��?c8d����J?5�C�|a"�Ti599%�-A�S�����
�������@�_@�0a�y��o��t���2�2����c�]ED�6C!th_]&$��Wdm욨���4����T�+#﬜;�h�W�!O�����G��#ۊ�pĈNu�|�U���)YÇ.<��yĮ��%
d�� 7�N9z"����z�z�t�e�zx�\��o�ckc&����>�����I�,}��5���ۋ�e���q��}��Q�r<1ƻX}��9�.��l|6D�*�����������	�S�D+�co�O�K���s�;��#��ZCAP��b@�9"�G��H߰m��*؍�L;��7��R�HHC���(�f|�I��_']��Mݎ:;@Гc�uFp��U�+~��p!&�ˆw�dœnt���wK[�.�@"5;���!�B\�k��p���"�p@c��OĄ�[��2�����b\��h�2o{��:�����\���'���i���N��6o��%�����w31� �-j��\� ��EM�r���L^s���L�W��WtI�Z��6�Ϻ�܀�E�,	���1�Dy�s[7�+�!�����`ߥ�~���Jzso;�d��3zw�$8��؎�]�aR��״�)H��097�M��9I���Rb��P%�a���u�$�2�E��N�-��+���������f7��JB�WG)Ւ�0������!���Yk9rdU�ջ� ;�45���7���Kl|����x�����\���q����kwgL�.~v���-;���h��7���STSM�UAc�>O:Ր����L��H���Iv7�����������w0����$hFX�C!������m����m5��]�Q�Ze���7ϋH���m<��H��s��D�߫U	#�o8h�����:#_�ؐ��Zc����I|�#��=�W֛�3�9��`���sQ��Xn����Y�����.&��e�(�xP<�*�◠�;�	�u�5���=C����)1�P���I�&�oA�Y?%�H�F�s	iV��{���`z��< �/�K �w����� �'���6��v(�W4NPÝPAY��7ԵL��9��7��8?� ��}c,��N/���y�@~&�,����I+^��b��S�������=\%>�~�&#�`ւ�X(��`�yCB�l��5u�r���p��\���8��;�˗Y��ZtX�ba��h�g3CC�t�8�`�����2��{j�<m����
�O'��p��`�R���*2���'22�}�8���� G���.t�؈G0�D���-;s�..c(pڈ��t�h���gq:5�i�/<a_�@����&���N�0-��-�q��fm�fX:�v��c.�i��H�N^Q����R�:D��P�9؟˓G��f��dZ]�L,�VR������J򋏶{j���|��GG�[*j!�Gl����*l:#��SG	�Ub�cy$MF�B�D����dd�!7�R�>��N"6З`v<	��)EN�3��u7� u�B���`�d\�O�Mf�k�qCc�N�In;gIQ��&�e��0'xa7?�%I�+"� ��Fg_�S~��Q~U�G��ꭰq4�	��pB�S9ŗM
 �md2g�:H̉� �����������h�,�ɑ��9��<�F�7�����ܝ@r�Ħ�'�}���Ł-�6��'d��oz]��9Ί�Y���/��0��e^t�c�����f_J 0�l�@kJDw�i,��UW����D;($�4X���M�X�8�+���$��ݘ���3�:�ftU�Z��R����G�+��h��q���;�=�T!�mJ9Q�����k�1��V�j��~�qX/�	���,�2nr���ġy���qO*C�h�?t�����H_�uØ�@�)4�;N
�B.ǋ_eh���<x��>��\��y�'��3�m<[TL�s�z�:�uG;M����������]G��Xyn2�vl��zcxJ��K����	!�٦\*ٽoBK�8
R��6��<�i�D�h�Ⴡ/��F橩W4�]���'-;��eo7�P[�j̓�mr�o����⅛��L��������6Cq�d�K�P�#��/	b������T��v�@|�{-Rt�ۓ��o8�J�����,�Т�Ϲm=(-�8����Ԇ���B׳����N]�ލ�_}�#�Tt�֛�������U�qh���Q��QIO����
����Ei&4���Z��i�d#SWjRDz����Qv����*[6-���w^lJ{���P7���t�_����u���H] c�"�,-R��!V�[�>���m4��&W:�����F��u��i�i���� �ӝ��T�zeM�����o%������D[������!�'�O��v��mt�[�>��ۯ��(ĆF�L��b4?߀3KtQ�f	��ՑG�n��64;�*L�����"{���B�) ��X�V��	�#7����@�b���| ���A�6 �	։��|��~�o��x���`7k�{���J��.�Ɍ6��1#_�I=��i��B�H��g4;��D28��ΈV������!TH�.?ݟ"[�*��,�$9Qn�EVBv����Gb�nD�>NBx��K>��I18i���D����u]H��M;p��*�@!ղ��?�G@�����EwB�{�*��ϯ��F���W��o���{�zm<y������H��@���깶�����j�ͯ��C��J�ٹ�&�dCaJ*��9�@n$S|V��;�N�Wj��:Hk��Z����c��������ϣ�mc&� p���f����!��GiR�cY1�JaO��A�����&sl��ݶ 3&���Z
��|2������ �܃k�䔭Ԧ�/&+뒰�E�T�9��<7'�dV}��� (�����Ŷp?&����F�ߟR4��%��C���(�WmS;�m�}�$N�0e��U9qLԖ>�Xn���2����)�6�ߒI�v�e`�t��v �?���l�@=�gX��-]H8���{�.�i0�m���t�Q�W�k��3.(��>>?�~�}=�~��BS�44j�B���<!�Uמ�6B��:X���@A���Ӵ��>����^�ȦﻡB� dQ�7_a>6d~�@�P�aP��u�96q1k��z��Wl��dE"�&1nmuܵ��H.:{������q'����5:��2C� ����c<b�%(�PB�:�6�2��е����OQ2fҦ�6X�-�`�s���g��^�$K�뭮L1���T:��z��MLpnl��p�$jn�y�f�#q�b��}n�d��+�;���U�k�?@���t�Q�"�l]V2\�֧9l��@������_���y��Ԙ���z|���`燑�V-U0[��۱G�7A�A.A{d����ɷpzۃ4����y��B�����k�,A��B?�������5��R?_����D��4�A笵���o\�@�
*7�������������r���ܩ'�F�CT�Zv��|�}�uF����w�V�m��/1�ACo>�ѕ�-WG��E��~u<�<谑{�	8���. i�m	��ƈy'��}���ۂ&�z��,��������pxg����U'7g!R��[Ed�V��@��c�'Ę�z/^�<�,�|u�`��� �#P(3d�xQ���1<�k%����HT@p޹��n\l���?��SWB����_�O~E���<��D?���0(�.��-������h�Z����+���/��.���IkL���N�@iu�En6صw�g�6Z���.��j�s�C
z�n0K����	�c��j�Ì! '9��s���H �#a�L|�Z{��<�5"(�a��5x�0�]�����#����0�t���4ծ/��S'뻫(�j�&'�'5�Ne��1]`B4�e$>\J=��5�D,���$��l�5����Z
���K��p�1&`�������������7~�Ɇs��X�y��
���Ы����3���u@�̹z�u ��0��R�r���r�VӺCf�"��LY-�5�N	�G�S�W<ڭd���Q���Z18��#���2;Ȩ��of��d\���`:$�^`�=.$9�7C=֔n�~�I:�,F���Ђ�Q�M�u(��������Y���|�C�n���-ĭ�%]����l͆v��[��K�JZ?{�K�^/�[�g���	�����0�kgǟR�.� 4!��Et�U���@r�%��`�$	5d{�3����
���[�F��M�G������N��|C��f6]�wp��W���ZynndG;�]p��ӕ�'��I:W.�a�����i�f� ��m��O�u֗@],k�k�A,�gn�9X\����j�j��mռO�rz�5�сG:��X����Ө3T4���I��:?@cx/T���.�/���3�085)í���� &@�L�������bZӸ5(��5�l�@Og���5�	ˋE0l��O�c6�K0;���-t����|7'w1�Gn���E-C���ʡםSBc��'�k�.�\�;�p깝����9b�j_���mʶ�(��������c.�In!f��7�A�<�`�^@��O�#b������A��`Bw��I#�9
OV-�NH�������;`�r�fh�%�'�<���K1HQ�W��+v����9���/V��#*'dI?�?��R��޶f,��#��{Kpd_*��@��!��f:6@���	:w��Yq�o^-J��k�B��{��`f�!�Vq\Y��O�z��v�{>zT�p��ɩ�#$Z�p�P�e<��u��(f��-��	 �{	�>D���^�m�3�c��%�'�ÿ�+��%��a�fv �"�M]NV佄� ��_������R��ܚ�mv�m52�{��-T�:�,| &(�AW���(�i��;���Ky 'W��������  �x]�
��k����|f����ޑ��Ib'x��Ft|���f��Ɣ��V��A�R߁e?���,�;���$�+��`� 
����y�d�BRv&���-2���p���3] f�VJN����؊�%6��NV�1��[en<8�l���!�s���+6�6�F�D`�
/P8oভۥ��V���E������R�e��'��e�v�D����9�9�|v+U�/�bt/@�9%�`J�L윛	Zl��g��T%rG��� �@��辽���$)ڲ�������8^Y�j���q����k9������*�A�
����(�\C�Wʰ�|�]�iZ�_�T�X��pcc��
CVf��G�:�dZ&���>�W"$��\A!n�S2y�Y2�PK[K"T��S�u���0wK���<�	�����﹓6(���{��y�u�5a���Vx��BS#��I���͝�.z�h�3<ρԽ��m贾�I??'dZz�X�F��O�^���j�q�;�=
f�L�F�H	�{�.F0I��g)e��J�Ş��;���\��O�4b7P:�����qY�g<���W�V� <��O�N	*�M�%��*�e�Bث�G����$�T���ylTA�~�K�T�R���^�iz~;���1%?�3Q$����y��qUO�2hy�ha�fw���c�.�����si������ 1��F���˹�l7�+�~rr�7菓
NmwB��沗f�MH7E���O� ���.Ĩxh?�]�y�c&Rn�[�v�.�	o�6ƈd�:�����Z��|��B�bM��J�u�C�)�G#�"j�E�d��"��`M��a�-�锫2�����EW���5��YRq�㛙<�/���u�"��W][&��/gW]w�`/J�P�|�1��N9��
\k(������JuK�[*�n�&�ș��uh���@� K�^�E!p�F�#�ː�t�Jc�K]+Ǝ���,?��1+��VQ�-emEp�a��:ENz1��9C= ��	�:��K��nƽoN�{�g��0(�-����N���N�:�4�͞��Aqן� ������N:�z��K�y&�����^�$�!��G�Ԡ�����D���;��2xˏ�s���N��7fh9��D�� �@5�ڑ��PPC-��3C����F��{�S�I'S�L�JY�?��G������'� �M՘;���������P|w�rCN�I
�J-��ODDB�T�n=��}�%B��Y���fa��a{�o��`�p��f�43�N�
wKpŷ��4��Q���a��N���@�nM�[І�{���_z?Oumk��|#�����J��@x��ŊլU���d�H�tC��u��'	؄�wD��r��q�Z��1��F�;�u����{*������"��[���ء�Fa�֛*\�����u�-�>>��N6 Js&VD�!�GR-��]{�|�r���@��y㐀�[���?�9гpB���E�@rOUݽ�����i
�PFL��8}���Bz�شI�^<K��aBvd����0�Ղ���U\�?���mW`��0�9�� ��W�k$�K��K& �p�Uo-������ǰF02o����L��܅���v���H�lg��We��*��nH=��p��wb֤:���a�מ�M;�w�l�C��o��3�)[�85��������;BUߛ|]��Dp��o�����k!�~�Nj����V;������s�
��<��{τ�j�ϙ�_��dw ���=�S��X���_V��'d�)܃�pJ�O��0g�2Q�]�n٩c���,F��^�s/L,"�T�'B�4�B՘��Xsm��;�v/ ���Ο����d�H���$�pfWb���k��U�j�>u�ў`7!++��%��~U놴��xn�Wu�����4w�/��E^��!����1�8e�o�Ҵ.�Z���Q�ث��*x�g >(v�1"���Vc5���,�V+GQf��~�b��'�:L"�-�ji�~��7r��B=T�1{���|���66��.���.��?�Rĩsy^��O�M��_�� nDp{Jr�E�V���͝���_@k���Ǣd�8m�j�(B�cn�"tnkV� Es�q{���ʂ��{[ڭ��4�!XcX���tb�eo�����v=O=��!=���$�(�i2#p�˷9wa�/tk���Y�>݋	K����J��ʋ΂��g��,഻C��\x�{�]�3�:��F<88w%:��Bϐ!�1��rD;Z��=�k�Ñ�����}�4:��8�Ek�*Ʉ!�yU$x�+�.4ͫ���I5ڞ PlX�H���`�W�m���7�[ƺ\E��s��z�-&������_�0���uMSS��X�HWBD�CL�������L�>�ea-涞��'?v��S�g�A�c��K���e��ʊ���r�>'H�tg�`e��]���ts���~��S��JXj�f����f)�}�_���G���ʟQgVh�<ui�5�0dB�#���U?F�Ĩ=��<ky�!a�Ti�ʻbdwR�����;>�-p�ћs)|��$���N�/ �QŝM���H��΍a�9�����Ұg�vL���+�   �O�F�$@Mrʞ�??;)����[b�_�P�h%�/ٖ�������c"��h�A�v|������rJn/�~<[S"h�%��Z���
M�"e�Sf��u�E��'��,~��}�����+��pWB��v�m�E�A���Rv3�D�`�H#�mQO��s���*g�B���'��~��i��Ů�)���Йꘊja�Z����Q@�$~���	*��|���̵��iR����)l��{��!�����M��Û�+�i@^]}0{˾T@X�^�?/��Y@��{�����f�a"���HC�Rɼ�͇B���_�Q��r�"������b�|�����b�=�O6Kk��*�M�g���/���Xboa�s[1�i��2�_e����f9f r�L�Ѷ�uy��lt���=|�.�ѹ�.+�� �pBRh���^��`:�)Ȋ���1�����Y|[�c��F^��9:9m�<ˇ��(\�M�߈f=�O��ΆF����}N10Hgs���y�T�:�eYuS��_�,�[l���T����"��G�����)�!p�s1��?�&���z�� ӈ�X��	�^�3�J���	]���|��љQ�M�E���]���A��<*'�R��]K�}@_���δ���S>N�D�i�L���(�g7�c¢���[��RL9&0��c� ����$U���%�n����]�[�4�=��{V2���.�F���4_m��nѮ��J1�󖈆d顛�N}k�⮟ �^ �扅U4�9ɢ(��O��`f�����ĥE��^7O'��"�PAp�U�(sL&GM ���33@�_N�ۙ�����E-�W�g|���B`.<k鳼X��5[��ș��h�c�y� h��7r�:��>:�H��>'�V��U�,o��T;p�7����CxL���h�H�s��z �3!���?����q���� ����/B��b{fx�Rt*�����ɇN����N|p����(e��]O�_X�Sn>p�z��D.�@4qڗw��#S�y�(B�n^,�?�xT��i�97O�/	1V��Y ��)�ՠUe}^�'�d���o�ؓ~Xfs��-u�^�0�o�[/+$�ŭ����{{m��������~8��j�
��Ƌk�Ƈշ2�M��|���l��D�	_|��7YV��E�����%�"�6�x�@qBE�� Zwd��>�,���������=d��I�"8��͋�,2�m��2q%���p�$hd&���I��f7��lX�lU�O<w�a2ـtǉ���l`]����c�g�}?#/:���T����b6�]7�'t��qG��=���b��R詔iDY�tP�?��EkA"~���3�u�<� Y���Ƀ�x�})>��
�Ƿ7���Z���+}�X"�P+�$���}�����)��,�R_�Vp&(o�𛧍v_Y*�����f�����r����Q�������}�q�o��7�o ?y 7�r����^�uf���ċ��V���� �K_F�2gO�Kڸ@S��ε�<���/�x����^���uUW*7�0��:eq���\����?Vl��֚AZ;�� 2_��!�٫�2�e��G�8��ݤ;T����cB=�L���&e���1�Du�(�����D��å<oފ�Z�����0�`�N涆^�1�y\��.���aEb���5�`���u0�������C=5�&�c70�x~�F$ Z��^ #/
wN�bȻDJV B]k����'�U�Ǖ�?�@�ϋ�]��5��Y�i5������ω�$@n��Wy}(L�V�d�6����f'�%^,�yEo�v�;���i�|ڟr	I�:�mbB� ��N���o����V�&B�i��Ὕ_Ι8^ϭ5Yy��]�u_Ϗ-o�<+�V-~`�u����=��k�����j!��-j����NX3>K�RMr��I_p���\dܣ�E�O�E
����s2yg |W9;�z&L`
<�wiF3�d�����U��6����dG��p��ǟQ�d�~�Ǟjz��]G{��c�	=/�mgjq9#����H��Zm�ǹ4�;�O����<u7钔�>S�G������t"ɑ�1p	�Q��G0�@�rE��_	�֫�b[����w�/��'x��}���.�7	%�ߒD[�Gڷ*;����7�uoA��|&xxv>I(۬�C��D{��q�MJscE��0f k`�c{�o��sno�M�j�>�n��>�%�hpVtԚO��I�7�$�1}0¢Av�6���NE� ���W�^��SȀ�P�-������m���'L|yX��a�AOi���p���s�%��(��X�I���@�̻#~��-�f�a��=�׵���zq�G�ID3�wB��/�J�p{L�M�Cߖ��>%�N=�����;����؉I�5e[=k=^��;lrxx�*K/S},��Al�Sbc�R��r.��� ӳ8/se�S�J�'H7J���������U����Y+���Mj���oń�:��+�u�{=p���'�ӫ ivLPV�/�?�
~���kr�L�̱k��i�y�?�9�8��x+��jt��2�D���$��%��*�/�zn�R�
�H}�`�9���o~c�&