��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ`T�}�w7�ɴ��劂�[���U*i�:����T��|{*�F�E�Q��d����3�6�:r`�w�O�oEޠ�9gr�8Z(�V�7�Z���W>�����TG(��t��qs���sb�b�Z�)O@�5m�1��2\�Qg7���|A�6rظ����N-@	�g�9a�y{�J
���&K|�x巌�S��� �Ƴ|��/���;�֊�}],�(b�d�%���z}�;Ԇ鍔�=L�L�i�O��&$[�����c)>3*>�B-W��D���E��{�	6�2@�[5
����>�|d����M�o>�򑍗�a ����3?-bk��d�u%^�=�<��U�]S�(}�Q�ѷ%��GOh^`�e���NvJ�f��Dt�m'5 X��I �Rh��� �wM���n��f�<�(������e�,&E�����0�S���*��Ĉ[�ߒ4Cn���t�M�w�,�z�ޅ�WR�x��Z�������3��H��0�eC��O�a��ԟ�|3lT��$ ,��������7�tR��c?���,����&[�2��HTu�3Q�ݷ�c�+d��ۥh3Q�F7��(�ڃ}�3J=B�F(�Zf+��"�q@B$t`'���r��dTFjg?�n��D�����vc�A~]��AXhh�#p3/X���������Gn'���h:�p
+/�N ���T�ց;ե����I��>�E0�c�D-�*����\��a�,��H�q�aӽ���#5��ju�F��c�ᥥP%��w�QE0��Bh��!��
��7p����}���Y8��1��QSA�l����V��Ǉ�A�>`k5���V�Qpn`5.E�H���՜���>�;��݂2@K��pb��+���'XWuh?�)f/�,����*f/,R�����x�� �R���+Z'�U���+ю�522YR�fM5����W�}�V_8$��~4��@>��1��ʡ���:��#Wq�o�4�8"�'m`����O�/�+�6�m���t˿k�\i�# \�/U�p����׮_C�@#)�԰.l!���N����8�Z����f��ǧoY��z��7�Ǯ�ӛdz���	�� ��=�z�P���í!�1l�zR��,�����j����x���J�=�9����8��ud�٦)7�Q��K@q�	��GuO\M߸�S�vq.ݕ	�8�T��@�4��H�]�),՗s� MO������g�`�Lf�d":"J�X�$O-s�,i�P�?H��7����D!�xR�w���(�����D����dkqHpq�{��$QntY�n=��^���ў�Iu-	0�x��m���N@nB8~��O����z�����-p��[�f��>�'�'+�i��z7^}�J"wXNJ���o:���������v˺�9��jP��u���v`�?�8Þ�"-�����f�m&��̴��I�YL����ia1-�Jh-ZB�[#��Zz�/|��b�(q���{��gh�[o�(]�� Q�ȢJGM�]6 O��C�E;�۷vc�~p:(�r*���C��
�dr�����B�5!xӷ��ߌ�`�#�$@}��K����,3�L�����Û)Hfp�:i��'c=���(d' ��}aԖ߸C�~�H�Z�}loɘ��� :�����d�% �G	!)ႊ��6��Es+��U5����/#7�&p	����z��ɐ��<������ugj؍8x��a%�|�y�i"�\Wze��y�r/t"���j}�����
X��"���GD�gU��P=�$ʲk�����I��"y�.�3.�i����Q������X���D�O���uo���/t�;&4�Y�.��bF�܋�ȖOSQ-)Y�>8ʓ��V������.��M�T<�;>�2��M
�y��*ڔ�v��Y�T}�xzj��1oR�H�PѢu��� �mo$�}�H%&U�?;�����<Q% �u\F�V�k����
����~����e�x�ǦEsog�c�8�W�B��SP005������en��jq:�J���w�|�>g"B�rP���������<\3]?Ţ��0�5��5r�����Y��/JIYti'z͋����~���%M2s�we��\��.�	��R���'��F�c}����Ūݤv2ו_�F��v�!f^e�?�vc�1�jX��"��'h�%���3_Ω�v�$L�*�1�zG^Yd:{��'P�Y�:!����ٗS><,�n����Z�!�C�{'��p��
$�X��H���*����+�<ү��/���\�-�=q��1��L��	�!�+���� ����ʚ�WѩS�kkډ-��1-/9O�*H�Ѕ�����%�@�x%�Q�?�z�%ظ]Z�)s�O���h ��Ps��L�����
K���:~s�<�u���t�	Z���5'�s��8��<�O�%r$OC�B���G��T
��;|u+�3�ګzf0�0!�7��I�0�Z!�N�G9�εY����d�@A��좧�-�q��4���!�RE��>r0�c����V�$�XSы����@ �;�_�`�x�1W�������`����Z�:�2ˡ&�x�+��Z֩WA��l��E�{��E�Q[��;�1�_=���X���$hmS5	��=�׌*E�����H����\=�����l^����9�	t�j�GXc0Gaؿ[݌.M�����t1��K7�w�����%Ɩ��4W�R���'�l+rH��L�Z�j�W<�	�CI����cS�)Pz��䉒e��p�ۄ�w>Q%*Gc�ʰ�W���3����V��ķ���d��c�dؠ�p@�A➴η0	7*nu��h��pҺ���[^� t: M�G�ѫ��{���i"#�T���g����9�"n:ҀU-�jLìb���,�:�e~��T_F�Hn��B��C�!�bj��ő�?*�#u^�g��gۇ���c߈�=��s�۰K9����2�5p�8��#�;���'�F\����5ȄXl�>�Q�i>.ͫ��^��KF�omǗ������v����ْ
��.�T��9a�/O@���{�X@X�K��D�U���W�F
@7`L�#S���$����_�u���Η���-�Ew>�H6_6��s'�v�޿�#bfv~xf78u�Ɣ%f� ���K�#T<��/��6���V"x"Axc�T��j��D���Z�e�᮶�x�M(�/��-U���1�"�⬿�(}qq'���x�$"Ӑ���=0Z1E�i\�z��,P5O7��gB��GQʦe�Y-�hYu&9����tWr찙m�� ��ve�
Ց��=�g�l�Q&�@_��=������m[�p�R�Ѭ�uБb�2O��*5+n��a�\J���﹜B����=��{�-�a2���/���Ǫ�!���UdF���}�����l�_�������|��O�������ܤ���s!ŉm˄��'O.T[�|�ùd��a@q�6��f�y"��A&���P$G����qy(Ƌ{�􏵼�P��C�ˀ{
i�l���^FQ��w :A06~�q\�'g�N��J�D�v1hzD����\e�| ��vX!��'�-�j����0��@V��?�����#IB�6��?=|�-���F���'}�2�ٖ��"7����h�d��r/ ��mK6�t!�<�]>��U�.����xO�_�K�5���t40�0�,":�ʷ�8O�[���<���YZ������;�T.
?�_�=�V�Rj��d��P����F�Ku(��&��Y����D��c���4A;��˝(\�Ɏ%vP����O-W���r�����7Ӄi�A���:�)���[�`O�74tRWq>ԣ��3��B����r���n��>�Y{���)�| 5CY���x�W,�����9����iVhkg(���b?'_��_V{Y������/��v�/T�4���͉1����,%@�O���ݻ����Hث���8�����У+F�{[��� Ϣ�F�,0NK���G�N2��p�.n�<�+\�� s�11ߧ�q�?@l�n�{\�Ҧ��VX�d�Z���+�Ə������a��%_R���\6��#�ݺ!��X�Z�/��� 5|d֌��ڊn.�9�Y�k¸����M��D�Vu_{�g��)�qD}WCO%c����坺>B%�~@4l{��}��ل	p���:�`��t%$��.꽺�y���S�Ȥ�+l��0	}�E�)ɥaHR#R�j�2/�4���K�i�e
�gw�v��lP(��e\�n|����o9h�M�k�z�(�K_�>�¦�>���=�(��/��r�t4t����{����3���P�$9�^6o��oV��>dS������lH�#)<�'!r!�oP���,�w!X#k�.�_��b���-[�0n�P"<�Hk0(^Ӧ1����[����:����$3 fU竈�F�T�u&�
c7֯k��^��WnB��1v��c��z��Q|�%l����P�Z6)���	h��WÕ~�_�P ����B*=`��ìk����¹tĘ�zf?c�h;�˟B�%�#����TT��W7��	�L�~Z�r�����j��Cxq������3�j��Ho��b*�2���~�҃Y)y�`M���g�|y2�Lˑ�4�L�.��Q;�=s��W5&��U)�6<�B�P��6���`�ͦ�;t���Qڨ< �.0�.�"��E�&��؜��:L�����C���8<�39��b�o%I�p�Mё,o���7��%�є^�q����U$��5�ʑ)Hg�ǽ�A�K�hH=a�eNh�\H��x�����g�Վ��	��"<��C��R'�h������q��HJ[�����g�)f���w���k)�|���4�5|���	Y�e ���p��E�x��X7���@��]0�_[�����f��\b�@(oCнm
��5�@~.���+�FJ9n�޻9rm<�D���ݮtrh��Ȩnu���Ȇ��:헠�Q��_s�+� �S5^�n�H�y�n·� ZG�*�*6 ԍu�%�}d4�\%��?�5��'��z�u��O$��鎛�ʮU���7��p#��ڻ!sO*�|NQ�@�A�E��Q��`�:L,���@6��To��`�����z�����_Qewi@cz�y�'M���=��<�/��8ɮ�y͌�D{�!��&	�=�6�5|J�n~��5=و�/|	�H[t�Z�n:)��s�a�od�YV�G�U�cǺ�m��22�� �.��oem':���%��`�<v�17��Mj�U�O��3�PF�1d�a�-��>�Ѝ dLK�I�ؒ��E���\���[��YѮs�����Y���c5�S�mb��?r��|;"^��C�+�氘$��)��1=e=h����>W���IA��^>���u�Y^8���9O �r�����n�N���<����i����
!@��t��.������)��u��q}�d>7�gѯ�ر����If�y�����ܰ���Ɂ��x�h�y�9�c`��B��	��&���U̒T2�`�tzK�:lB��1���_��I�T��L����O�D@J���X�����7�Ya8�I����6���0�oy#^f������T�	�b#=���p`��0B�k��G����ݨ�9SF_o�a
)�0*&a�{�J>0l<�z-���Q<�3��ۅl<`�.��$Zu�H
��3�t�">e���ֶ�\�1	Q��94�p?ʙ������f��=���d�4tpq���M婐�h�ˬ)dyG�9�v5��\6фN��m,C#�����rIo�LN�u��s�� g��ƅU�i��-�/1[���C����H�~��2����JP!봮�웠� :��3Ɩ��
i�l �7�EO��J����\��_�;Kh-k;����!��:#Pr�ɰ���fMo4��Iߑ�Q��d�
LT�cJ��|m�GISPh�S���/�>�1E>w�k�֨`�����ej��;�	X�M��%Ӆ�,��������~�+�=�+�4�V�r��m�:��Û���ô�B� �5�k���5,���H�)�{($%Vt�a�������γ��:j�`!ߔ�!PM���6j5RD��%&J���/�ݢ먗�w�IH��oCdz�a0�ٗl��mP�h�:lbu*[S9sgֶ��D�.e,$���\���#j���D���FK�o�5�vs�^��j8�� �yi��F���@�{��ۜ0s�t���\KPႚ��$:MT����N�'x92&���{&L�L�Q��[�<���X�S�����.Jv�N��>����]-�
�l��8K�ޚ��;+pM�>j�*#���u1=�7$p��Kֺ�*ʹ��@�Z��q�jvW�5d=5e��¦U�������_��N�R��՜A1xx+�h�1R��E����2�/r���P�������Ջ�)qcj�}0�7�Cw�<�O�,U\�k���l���g�\cC&̲'kd��[S�����J�遡�'?���U�J�F}�j������ӚU��4d��%���)2G��z�D�/�*';��+ ˮ�3�L���-!�����[����D:{�P�j��Z C���-�Nb���}�N�$r���m�֣h}��.���H�5NO�-���8 fÅ�IN�{�����呏���檿��� �+�N���/���',�mY���7�MC��S�A��s�-c=�l��ʝS+N܃v�X˗k�;�޷�Z�f�<X�7�r�������a;5�=�9�}�%h>\������~����g���|�w�x����0&(�)�1�7��f�jQ�+��B�V��w,B�c����V)[�eF�c�X@�u��v��lr�2��j0룁�J]���}�A�Ր��6c�����5�xQ:�iز��2���t���e�$��+⏈�dE-?�6gS�r*��\�ې�o��5�e:�(u�D�S;����/�bZK)���i|͎�}�`���*A�Jr;COiG�/J�Ź �}�3�l�����<_��VZte��ޮw
\��{䧏�v�R.�����QM�S�`e���"��U����ݻ�;n�m�b����m�Lİ�O̥��� B�VƐG+J"Vx?�%@���ݭ�����x4w�Op�*��҃_�W�.��y��ZA?�\S����N� Ku֊��
8f�N�	,��c(�e�K��(��k�ei��L��&K����С
o����l�&݉�d�L�8xG�m�!���@��>��u 7����C��}�b�)=vY��ӊd�R;��[�8}�]`�d;<�hB�Sb���/����3��&g������|�������p�C��'A�4l#D���'��Q�304�.����~�`M������r���x�y��~ah�)�q��HMܡ�y���j.����8��Tl�<�Bh�O_^��qN�Ra����р��������|:���ػKm��HO��� ?�_��n�s-mK����{zE�l�u�u��E��2�͂-)a�,`x�R6�� v8M��St(`��Jo��N��8%�A�zL϶q%����U�n
J9N�� ��*���P#�"��b�&𥩃�ӎ�P�����ع�4O�X	 �v�'�����zs���~^�(SU�e*��Usؿ��y�9�H3'O�/�Ǧ��\�R��Г��W:�|��s���
�>=s!�/ d�+"�V������"O7��\k)����>�:-�A�᫤;�Rt��1;�<t���o���]߀Uњ�b���t��?�MNU�UB��r��t�yK3��QC��;W�2o�͡�[,�M���H�ˁ"����S��p �ܒ�Qd��}��u�P;�Hu��e����l�����fgs �[O\��۩_%x!y��s`�h@6�K�p�8�����T��ߗ�Nw�����d}63��U��XϞ��T��Wt�@(vSm�)c\*.�Yw���'d���q�c���J�;�_��e��E;�Z2"�����2Z��!ǩ/I����*���*p�L�<���}w]��|S,;M�^��� ���j����pU��5I�>��Ϩp�N�B�	 ��af�'��W�kÖ����Cj�{��%�����бU��To�|NՋ�×9�{�E?�����:e��z�Y�Ģ:cj)�KGXS���O�].���ր]S#�M���d{Q�����<r�k��K�C%2:YߛXI4�O
����TP��Ls���m�FK�߆xŀj�fF�̥��/3���c�o?$�>P����ma]�ܔ��X�߰Q����#��&޶z���=m?��8
]`}3
O#A��za�%�p<��b=r�����~�I��ZL��~�Xgh�F&��t�S�ݥJ������Cg�J��+�J5`g�pA�X>�t��DN���b���A���G�	�bdi��_�)/�Լ��\r�Ծ��q:\���t<`ẵi,���g�
�nߑ��U8��V��p�G5J@�xUKZf�!`f0-��9�֖%�)k���{�B�j��d�㈍ I��R"���1l� I�gK��`F�D���d"�S<3���n��f���qΑ~�=H8�m�>b�{���wo(�I���:CW͊�_�s[��C;
[��Q���(QI��
��c��K�<��:zr�/C���0Q��
P�_�J*�u�;�?�G�e��[�zqV�/R��c.޺~I?���
�!��  ��P���w�������s~0�\d��A�G�
�O��Vu�V ǉMw�)ӏ��Aj3������\VX��H�N�Dy��Y�h!&>�H^���r/�pf�j�R`��J豢g�-�&�bA���ւ�:B����jҵu���&��}�S�X�ssqa���u�=��ha�em�Q�@X
�F>�iC�-O�.�7:����zO�xM�֍QO��r'L��?w�ϐ�N��^� f�n�"�� ,w���;�4�������[���ԽI���W��eCs�B�W���ް*u�_���H���XP�@eJ�`@|�9�U�P�������:tE��̊����k�+�>N=ޢ����@7�9t-[��Pzf��5D����,A���n7��7���AJ�PMd�ۚZ�0����t5m	��Ϳ�bQ��aĘ�Et�^B�d0(�h�8�%pm�c�$�8��iSzWT��歛��\M�7����W��A��ѵ��V�O���h��L4��ی�p>,�鉢�
�G�]%�u�,��F�!��1ڽ:|��/�ʣJ���M"�$Ԯ>i`�ɽZy�V����{#�Q���eGN��+���� �\�ibX�~�q�� �v��m͂�t0�4".P?z�Ʃ�(n�%@2�l����1�qxз �]����6��0��C�M���t��C����/lj��v��'�a�:=C�c��N !�y�x>!�^)|�qP���m4��\:�6
�.fɹ�?g3�A�3tŷ�i~��b��n�P��6�3ʉ?�T��˵�=+B�+�8�_��' 40��K��
g_�kBqG��P
�L���
x�v�j���T
]o�|3��}��.G��A�=�VҺX~����m�m���"��;�dJKd�|�Ģ�-A~`�d!Ѧ�-!���<��h+#�q�!����E����E�$��Th�d�>�;(k�g
���p��5"��v�d"���R��pi2S(�o�eA���rH�J��3;.�*`A���L~��[�ׂ@�{Q,k��G�PӘ�<�{9GJ_B�Œ�'��@(_�Bv�-�ha�ڿ#Pe�례���J~���B������=N/]cu���'!J}�z�����d%i=��i)/��l�IN-�ė�=�qv�O�ލ�1]4׈%�$,��_I�?�����G�΂��>��
*u;��I�#�L���̋s�ɺ��vrXȮ�Z��� �იvnU)9]S��J|o!��B.Sn�$i����UV��kH��1d,�M���g�
�XU#�Q%����gϘ$7^D�2��L�.��V�MN��I����h+$�(P��X�>����8� ��>����Xl�"#�zGеY#����V��9�lǵ������Q�1>�����fo�s.t�Q��]AX*�Ҳ���~��=�y� �_���eW?�����0�M��Zv����"51��Y\�/�i��/��C�`�����+T�ܺ21u4��siq��Cj�faW��v[�U`�É#��+ٿ�]s��`�3��88��P<�'���Y�� Fd�	ޝ��ުt��7�
U�Y��h|���g��߳����|�$հY����+�/��1Ft����J�����i0qehF����ﺬt9��A���ct�T�KO|�7,�2V�H������w]]n��%�:�n7U��|��[�ǹśc���F>X���q���h�~D�z�xԶ+P-Y_h���ό����ҏ�e	��hX���7�Hߌ����v�*ٌ<m�
�3G��L��uL2����F�ȓ �w6�d�B �Ho�E����9�ZwRQ�� ����w��je{����H�Vǥ%^�;��B��U�Ef'd�n;>3��;�[k-�������������6c�dh��N�����r^&���BB�r0��:�TO 2�%�� :�B��Ȯ�U��0?��|8������7��R��C�x@b a&N�[T����W�Mn�x��܈��)�-D6j��u�D��#�S#��mBIvL� %6p�]v^S�v�C7v�YDZ�^KQ@��w���tht3`&� l�|i`��]����ICI��餰}DR�J���I/!�C%��i�,�}�ʈ_�:U-v���6�up��bG@?YL��_p�V7�'|~�5s����l;G��]���됎����?�c�
{H⾶��CaĞF�HvPlˋ��f���w����@��'X�TKdd�&,�����[yӫg�1n9��!���KJ������Z��1�A���%��c��zH��/[�Ͷ<�vF��p�I��W *����
�+�&���4f'��p��_�+ܼn�*�������B;��kT�>\�L�E;0��	j�c�G膬��h�(�8]5����ޒ�FM��H�Xw��)��OJ��W�돣��+P8�������Y�D�*}��w�0�ФG���Pb
�����B�4U��-Z �dQ{J��0gV`��֢%��+�癤��A<E����3��S;R>
1���3_d��1t�R ��wmY�1?��1�P��;��oT0��S��^���|YC����ʎd��v�֜�5C�Gc�6va>S���QԢ�,m>ƿ��!d�?T����W�&0}�IϪ��=8}�o&4��R5):�� iS+�j���|e��Wؗ�AJ_��$�D7}0�2��l�ɤV	s�s(�Ƚg���(_,�ѭd�j
�Ơ�`Q�By�d��<rd�I���&Uw�?���* ALW���U�D���$�;lnw��p[�L`��V������p�d�eՊ����Ҁ����l��V�^�D]��˖�O���Z^�612��$e��P�0'��1��3�&�
����t˶�}[V�ܽ�/+��W���O�GZ�d{��AD~���|�a����ý���7����1�5{n�w��kҴ������l$`j�.���a��޷-�'��N�O�K�a8m�ǩ%W����)v�O�i���.'�`bqsI "�n� ���q"�F��f�����N_����2�g�i���(RЎ�V���تBq3KJ�K��S(�G�8ǻ!o�N.����A���Q8��<6ᒌe[4N{D�����Z��l��a������#Y=�V�v�W�{�a��S�}��;�+M�g��̰��$Tx4!������xY29�zخ;�N�M�!��D����pC!>/���2`2���<E���`�|��ϔڔq�4��>e�ӯc�/�֍����q>gA�E��� ��Ǩ���
 %K.�8xm�\NL]Ɉ$��V�i�4�>�AZ!J:ln`Dʈ���c����A[��.)F�&���O��C�ۨ�KaU�=}^�O�ӏ3��� �]���N��:�n��W
U �7�u~w$����?pY�ʧ��`-R��bF�7�D�z1ۨ�;G���t�,J�Y�S�lIC5���)M����H0D-�fJB�V��ڌi�$���o�L��>�����Dn�6�Oi�3���	o��UH>yb�o%�}�i�
S�%�"�+��r墯n��w�ƅ�IԷr���yX��x�}g�|�P�J�>^�+ ����a�}dp
&�6"=���Ĺ�1���vm�����1iHĘ��2 d7��z�24��9 �Ne�24Ŝ5`��y����:�q���7哞��!�#�>�������e�5A����[m�K
F��ϐ�B��Q��<w��y�O�	M��ļ3&��Dt�JY1= Jn�{��W�~�@��A���=��E�'�9�B�2�U�V��5=11�"��2WOh��8��ɇ�6dK'0�C���C�H��m5���y}¨����eG�=%Y�v\������X��J�������Q�s~^�AV�SǸ��/Z�	T��hq��:\�>��9�D��ͺT����MB@2-�Zsȧ�_�k��2��f| ,eȦ��$�B�!�FcxL����ޯ�kXaj䔦��� ��_��V�P]5��F�'�W��aW���K�;��~�%bh̦�������~?4��3P6����d�QF�Ɯ'
�	���K��q�u��~捓{��N�=�Q�Hp��w@��b̬ }�n��z�U�
"[��m�6�E�� �}��ۧۏh�5[��~ʓ����Ц�Q㠰~;t�X�'���:�_G��� <���$����=��Qʀt�H3+h`C��S����䭼����Oݩ���㲀��(�=55!o�%i��{��Q"�z����+t$���}�ccKI3����|�Dr��<��
F*,��5�)|�pF m+����*8!��x�_��OJ(�����y�<�L���y�=��#79K!�+Z_is�O���t�m?]�#��N�s&����ݿ9.sų]�|C����NϽ��f�j���gКI���5,��IQ��`C�}�%2��	��{�"�b�_�z(�u�v�vΪu�`&�_ ����&(�mY��-��S瞙�G�Ju��]�����e��o�5�
@k᪷.%Oc���P����1W���id��{���b���]p
&8�w�g��]��b�@.�0�o�OYMen�4��<�To��]����P�,�P�pq�����fܡ�,ڃj�9w8U-�AM�}����g�ЂgH ���@K����(2$���f�� �'29uU�
k��/��U� ������:U��b;�;(46��v4��[J��r���|�C��8jb��8�'��|�S�����;=�P�x��x�*��^�)�
�Y�O�b�d��'Mo\B�c�N�+Kr�{I�����?'����Z�P�9єc�JK?����*}�9/�H�zIC�=�:e2�q�9�/�ҥO_g�Pl����DE��j�=���A�挶��H�9_�����B���]��b��[��� !N�J����} sC�.KIu6� M��в� ��
F�Z8�̤��ː<z���H�Ҵ��ٜa����6}z�*DV�,�h������Ø��~LSV�,=����g%�!Kc�'\H�
�_!�'�#�U�,<�o��"~�Ҭå	� o�.��͉#]���d7RkՍ���2�s�m)�c���E4�h'*#� ��U.:��)��h[,^��2��d��a#x�`�+#�y�+����<�.����iԓZ���v b�*��PI��,
�A���!�UzQ�4���8�9�o�y2�m��� IQ���x�h_:�_ϩ8�%�h�(�=�ȉ��[�1�<[��櫴�E�J���X����#t�`ur��q~≠HHz���O��l���8�R�r����yf��Zy��d���>R��V�<��3e��"�Wg����x}[T%<�AQ�V~Q��ˑ��'�����
�9������#�4��
!�{�hY�ĭ�`��sƿ���r#Щr��+&v;��)<�m���Հ�w �aI���5�v��sx�Y�=5������7f8�xk%מ��?��}5�5��v�9�����N ~֨����_��{7^��-oP�#�zԞ~�� &?V����^�� �0IL��*	7���ew�<ȓ��Q^�oYS?J �&ͦ��<�<Z��f�Y��im�(�����iI�w���W�"9	����������L g�7+�2����)y����kn1赭��ݼ��4�UT�HCV�V+��4$���x8�޳����&/JKu��7	�!s@B���S���TU�q2�3$���|9~c�K���R�fh��9�m���d&�W0S�P�����a��r
��6�e�����[�FG`*L�Y;�^�fR0���p!y9�pm��*$����(¢N��Y�F���j��ۣustJ7N���C����nj��o�u��S�O�+P�:��V�b��ڞ����̇�)�z�#d�?AF��j��lb��`���Oo��j�3�Ĩ����ϩⅨ�B��aA�*��tc�rQ#D���-�Q ��R��{�#~=��;b�5Z�F���*��ߒåf�b���M��E��g�(J�I��2�u�Y��d�ǿ:�]Q���ܴX8�8v�.Is�A�,h_���]"ȏ@$б�?�2s;�C)����@n��~g�a�fޔq k�F���
	�6�7}j�X�W�f�͞!�A����0�nQ˩�旼�"�;����1�3׶w�y�����BlƄH���3stU�� VK�^�_d� �a��������J���ܿ�^�kA��(	,G��/E͂AF��hW�0`���d���$MT$\��aN`�����h�Ml��w�F��Đ��{��;����:����֦�:Y���qe���9MU��Ɛ�ꊌ�sB�Ck�a��@�u����
jB*����j��-9��"ꆍ�mv3�-�~�n���GB �H�`�||�<��Rд����Ҙ�1� �@i)�wP�t���'�;��CGƿ~h�l��=�ďy ��Ac!�\Q�N�I�OX�:����u�7����4�}�T�Ʋ�>ܴ�g�F�m�����;V�^6�C)��A6�>�I�y~��_!xy6Li<]�����ϼf$=k+(�4D�D�c��4���T�0d�� �@)�Π�wC�G+�b�׷?��e��{��̔��B�	�T�ȗE�G��nCĺ��B��FL�l^�JC��1����`}���I8bc5��='Ҵy+ ���5:)�D�6�VD|حC�|��Lr�z�Rv�${��xD�˙ê�]����Q�h����q�*��B3�/.S����_��M�{��7骷J����(�%'<y��r�}F��x=b����s9�SVN�UMlSjʭّ��G�9q)Q'���Z�3�$�%�m!*8*�}@5�6O���I���3�s�y����A���7|��k,���x�r�B9{�rZ����\�T�s�tхCl� J�DfS��U�|A�V*6�s�=��,����c�_����[��1�c5���9��
3��S;�B�*�|�X.��5�FR��)��e��}=%�?����� a�O:v���KV����Z��;���o�I09��Y��D�Z�����4sx��A5���)T�&؅#F~���)���>f�u���{�ߣ�;���:�2J)����]٤��J�������LZpɪ{�V�exH����	��*�`ٰ�hA,S��%�U>H�<����(y��ZW��.��W�3n�J^�+�o���'4gh���?�r!;���ް=�գ7���V��GzK=�n�Z�,��оm0	����Ɋ���Ή����4�n1s�i��ٟ��	�n55������32�� �B���R{8F�T�Ӂ/k&�xhfS��G`�s@݁��V��&�m��\�/2�RijX^	x���C�>��E�ݧB4;�?�.6���hZ�4X�vժ�Q�S������˱��;>x���tV�̤hAq�tb�R�)���<'.�2�Kq�.A��"�6���b�<K�4��u!`�Y4E� �DW�u��� �o2	�TQ�S� %�K$ZFq)���\ᜆ��Fh��U���m�
��ʨ=B��\�y]���eIe ���D5����xP���js�~�1�=���F�>�Ы�o���]�.�f4��a�`;���95�`�'(��C��{�O� o�;���e��*��c;�G����(T�. =5p6���<1���Q�9�R��/+�"��׺���ύ�!���Xv�R�M�On��:�ۅ9�D	X�k�%���xZ!/�Nǣ�v�����"���7��߃P��Σ��梋h0s.�n�=|����j����6^��J�*}�Z5 �� K�er	�!�K�`�}�Ɂ �S�v9����^�gXU]�G♕!�����%zl���@�Bt
R*a S��٩��=�.�U�߱"�8\�^�� �%��:��M��ag>���M��-��Yϸ�[e�?m]r�	rJ}C"V�o�.��s��;��C޽(��BZ�l�dg{�9W⑨eD�쑼���NE�rr�y���jw�Fظ�~���`�<5���1l�e���IΜ����9)��jM2N.�)���Ie��l~�yO�v>V�zS��� ��bkhs������P�l!F����ϱ�����űR�3ۍ�l%Ms	�R�ĉ�E\~c4�2�d<�q���Jtn��O�N~р��#0��l���5�J�uF�t0��������/�Pz��:޼��̹��Iq�o�m����WV�$�lp}���d4�\R�
��
��F�k�����P�,3�6T5���Q�
 )o%�(�*�.T�/���w9�h�8��nP`������}��a�qD���z|�|��n�)�v%O�؁(��$��=��b�?��Um@���zwཬ���*=ڵ�0]r���k}�Be����/�׸7�w�M
�E�n�R����m��63�;���M�tY�dr�̌]���.}!�F���:4Jւ��j/���Q0�R>�g ��9�_L�_s&!Q�$����M�6̓���yt�F�|"�J���c鑟�#�����P�$"9?7��(\\�N������})�M�AҴ�>ԝ�7�Q��-[%�eWs�Jo���뗛wjU&�h����gk�tZy��{���?��ği.PCx�k��'}�{��@xr�,�^��Rڰ�ޛ��To6���~��c�w��$/��9T���72��eSv�H�"�Qd�Rpo@�Ʌ ��@�J�j���V�V:e�n�7`'0A��Spg?⑘���p�# b����Ǝl��'{�E����=y�ߝ?�x��-���B�dŢ:!!%���\	ո�7i_�UP}:0. �:��| �MbyM	�\��P_}=��]� @L�,����ح�X��R��8��0;0h���1�!���G �a��w'��ݚ�gA��c���$��>���u�!���O�M�Թ_�O�2��$���Y�-}WٮR�g���P���or׶-h���K�a1i�n\{�vx�n�;�W�dw�9����pRm����zR��i��uo8:�]l,\�-��O=
�<�Ns���Ȝ�3m�2J�؅�C� G
#���I�D�3�_��c��uQ�l��Vܣ��u&�7�;�̡��ir)v�Ҋ��gGC�\�1��`acL��N"DM�ڝ�u�7�їQ�& �=Mjƻ>k��r���vD�8aϾ$.$p�>,�y+9��n��>�\E^���z����X����O{!?��"u<zW�p[sֆ�]���&��B�y��@�Җ|+a�?�غ�
;+����/��8��y?u7���]�֔q�%^�K�����d��uS��Pff���w��w:���"���QFͶ�9e�/�3�\<�o���j�H��L��y��I�^\�Ny'����8�V����A�6B��˟)��Q
�-lQp���c�"�vK��y��`R��>��q���� ���A���'�C��7�?�xA�����M]��@J�S�����}�M���ۣ�yxl��2��1���N"��0G�=g�C�q�\����QRܔ������h?'9F��Q\MG�-^��
�AaslO"����Ua=*!����Į4�) ��&b�N�5���8����@�S��Fs;D�zh��|5O���C҄�#+7����L61�젓|(��-�sD������Y8U]�FcD�@~5?UWeC}p����H)�Ĭ�S/��.����W��C&��Td��!FY\�r�$$�
����<����7�Z�W(��7P�al�Y�:�h�t�xDY��T�?�����i�F�}���ȱ���[�&��M��!0��C�=Q�k��P���]�yU~�����b�&�� fZ�l�b�}sC��Q����y��p@��MpXP30����3�S�K�I��DTn����\��(%"m�R#C��QA��p��)�b���C7{��a�LGu�BR
� �b��	Z�uv�
�U�;��?wU�j���'���QwH�)��#�[���j���+��|I(gBRTQ�Wk�����r&�|8�#�b�����F��5N��Yv��n�����r��y�	y�;3��C�+���}̰��k�� ���8'�s=|��&�8!n +\�=��B2��Bod�	�� @����ȎQ�rQSs2�ۅΤ�S1��b���C�%��/��E�d���8X�gp���ݗd�9g����	q���a��"k��1X"xogY�{vzozwB�V�ǿ[VEI�ʶ��!���Ú��]��@��z
��§C��"�7��\fd����B��#��H���V�+Hf��H��4�g=u����k�M+���G�ê��8��
y�$��6+L�|����t�t�2�D�>q������	7���)JG��_�aZ�O�y�����qF��_�� ��z�a���-U�����,e�&Lo��� 19�U�N� ����GE��'�gW"[tc!��9ϔ�A�d�8s^�<��&�i}�$V?�Ď_�PCD	Bq�w��[���]��Y�������g�}�^�GΚB0a#��9(�n���M�t)��`�%9�<TBE�/�ު��.+f:���L��P�Zq���T�)L !��#&���=��p�A�Mikd�T��t[���čMţ��b�~�����S`V<��y�6��I�,Y�E|��w�[���l���k
;�h;g��Ѽ}"�Yܤ�D��A�-��솭U�	*����:<�:ݎZ�@��<ݴ�+�_5sYG��`����u�l�7�\Au����8�w�c��7�Ó9R`�.����7_�l�ӏ.��Tj�cj�J�,B���R��Kx��ր,H��hx������_��E��!�eR(GDS#$&a:Ė�v7��[�INU@�;���7��43�������!6�� ��.��1��a��6�*P��/n��9�;_
?�f�g��65�Z�+R}�����/dɿ./wH Τʊb�<���ܖ�5��2��(�N5�|s�P�k�"�Б�E&꿥�d �o��r{GPg��=�jG� T?��uϥ��'_Y��dG�w����5<w2�C�9F����%�'�?]:���"{�4���D��h;��Ww��c��WXXp��O�і�1�@$�紮�eC���OM'ǃ�x�F�L<P ��t�����r�DM ���܍W��`�&V��mK�Q:��J�%9�}�!�p�o$A�u�r��4������#� ��OWID�E�x6aO�C8����}���"b�d���>��(�UdF��l�w��������Ȳ#��u�L���?U6������.�@U
Sck���|+5iV~���::���$��߹(�hX���jZ��L��R���[3�-��<�rx4�зhcp )� �����k9�6N �4w5X\=���I��״YI�q'���IǑ��-j�Z�"�x��{��c��dx��g@���E'�z���`�K��X�����D�8J�b?HEs+{�o��0.��~�c5��ucBm^2?�.k�7�S��(ò$F	h7P;��%����� v�i.��ܢ��x[1[a'l\��'�?�C~s��;S��zC�ng� i�#��������B?�;<��8U�x,e�)�x�B���}"m�~�d�0§�� F�z���+���֢�3�1n�?k?s�<'�}_!��������dڶ�T�=��hX<b��%�z�w}m�����oE1�Pnz��2����FwN��5(~Իo�t�=�7��gWrV�3%�����5t�<'n���M��W�Z�`���b!�M;�X�Ȫ��[�+Ch{�F�1�
̻�X�/��e���q(�@��n�f!�y��Ka/#�� ̴+�)��H�� 3<��`<�|�zN�_��4){m\�F���g-@�� _J� V=��94A%�b,�'1+��>,>ГB�#����6Z4�.C�����`��1W}VsYޑ�.����w�ڳDet����`2��,�����_ ��wk)*k�|��GR�n�̣��� �M�-f����h�����$s�o$-�!��#��SV�Q8��HW���e]��G$Ef��K�@/#�s6� ^{�>��t��-Ό��d�� h�����z楏z2�WX�`�[�T�OT�̉��)�-��9�|�Lۦ8'�O������������A���D�$�Q�8յJ�[�����Áo�c_��T~@m�w̋}v��پ���D��w�z�K(q7���G,�Wb��\2�ݘ��9���G!x�3Kt�̎�}ޱ���a��p������ɀEy��V�^V�U�F'5*@󏢕�؅����t]���ݴ*�Gh�}��#���M�t1ZVנfkb�;>�+Wd��˫���f�ڙTD����4�(T������c�������������h��ş�p�,�":$X�3�9C><����K�M��f�bMݶ��4�~5�q~��)6�b!⌈�V`nZ����X�C�?tu�-v �P�Q��_�ȯѦ���S�k�'���v(X3k����p�{���OA���	Z�:�'ľ:f!��(�f��-
�k�К�"�ۦ�"ͬ\숔�$��`�#���I.S��� ��  L犬��9j��`�(������K�K��E����[��V�B��X�J�ޮ�2�������&M��Y��ͺ��>O�p�u��x����c�!}�.����p}��l��ks�`�s��-BCs�����w�VB*C�����m�J��"�,�K�ס�5b���+-��GZ,�����Yd�lF�*��m+�G�Ê�gq�И����+�ȻD��U�O6T��x��$��`�je
f)���W95�Ň���������Z��Ҵ>SP��HM�.Fۊ{�-l�ZC5�	�"r�uE��p�$��Uܰ��XPwɛ��Vu%ʷ����O�h��U�B�/-o��ٍ~�ͦ:K�O�^Z�����6SCd�@̦��,w��'���'S�툉�hV�2s#E��N��#]����*Q)ܨ��댘%j�\L$�,�qb��iZ`�6��b�>���+#3(��/!$�srPaDwl>���?;�� ���u�iz�it�͵Lo3!�\�߿����	$_Q��7��,�A���r+d�6��^(C�7�cɿ�)�<�㘮b6n�Μ����`-�j�2S���%3'�zD��ϼ�wL$�zFN���3+�{�'=�� ���H�����<."�M|]��HeP��ؾ�����g�4��T��`V\�(�|m���4c��%>�-��M,TBF�x(��D���8a^5�-���&^�r������g@��$|m����-�v�P�]v�׹F��)�ѫ�e�>���w�.��Z�谹_�� d��?A�]��}Z��|=��J_v��gE)�PO���yC�LU���-su�]{�
s��x6��'!&�jT��o�G��y���ثO��[�,y��'����è+������I�K��l�	Ԅ�!����H��	,zerRN��}�pL �S��ad��n�A�TɊO�jX���'ߘ�7�����/�2N�F����0�a,߃�I����	�C'���9�<̣M��ΐ͌��5WQ�!�6��py�y�Vq>:�DW.�g=_&�|e�@J�v��\���`���]�-^P����y��]�u4��6߰{�> Vl��K?em\C�IV�H���.B-7��>Q���W�-`�����L-��FAY�k�U;[o}'�1����,n�,duC����a�@}��:sBș�s�k;�oh3R�QbF��V�j�z^J�Z�չ*�CQ!u�)�~�r%ݴ��g@��y$����mkM4fs߆��\�~��Hl�r��l���b��\K];0����ut�D���*븖�'0�%�5��N����ξS�H�10;qh���q%G�sNa��9�^7���y�u�=�P�*+�o�$ӹ���`�����<�P��Ӊ���#�#�u�9w��U�z�Cj{%��.��
�r޳\sNN�� �O�V�����;@���X�#z!��Hd)M��`���Qز,/,��G+ebQ�[(�"���e�+�ݑ���`�l��}���ͪ=�Y���iR�Sr� �v�FI"@���BXB-�Q�˚1�>���~�U��iq�@S��(|�A�2�S-�����fM���N�L�d`��r��{����V���&S>>�����1�Q���6����+l�4�y���͏�	Jj���Ң����o��O.�G.; �x�YƱ��T��"a�b{'�cDo��q'%$�W)zF��TkHA� �</5��)�s�8���u�?7W�;�0�Ni�:Ԛ'�s��9�9nsz'3�<䳗���Uw�B��Y;I�5P{�R�3���Z������e����le �ky:��T���Z������	�>,J�r9зz�7'�����#��0~�_�2� �L1#���ʃQ5�N�b.�d�%�3�A_�<�P`�,�x�0�ml�����U���]���N�� �Wu8���3Ҏ�(1�x�߄͝�2i��#�,v�A�����ѿ���uh+�~ Ԏt����Ȍ/���h�>�W˽�:�k�.�ޣ�ՒE��+��F���Wv�rr.ب��-�� �e��b�~,��D�D�"���ہ��h�q��ҟ:qdv�����[����
�w�$�F0}�w��ٽ�0[��qa�7Hn���i���p�R"�N�0�IL���N=��Y-f��'{R����Fn=[ ������VnQ�rS�X��d�����Lr�]gJ|������y8t�a�%.m�d�c�C�������9U7��&�w��q��o�J���}=��?*�\͹�+�ݧ�B�	Εc���~�%'tN�����φ~���2iEc�<���!�Y��a"�-��MS�Q:��y]j$�IT�	Xɷ2�\|��0, <�_���7����zeZ�G�#k��B���i���#�´����%�zW�C����bF�Z썄�f�����I��ĎK��q$M52k�u�\sӫ;�unb���F�������-x��=[��c>D���. �I����E�7��I�y�R�{�39�v�o��i�1���P��������ax�C�iSH�2��wx-�.b���'�x8=k���*�AP0�)���"�N����n���~ ��n�Șj�4�Cحf�Y["���১i�յ:�z����D�����N�Y�Uvt'U���b0t �<�ڷ|q7���+4��!���N>!?���+��{�����X��{���Yvnz6j�5��O?�.�����m?�a�2�ɸ��q�ۼ|��߬�ۏ���'� -�w)݀g4/PY��z�n2�0��|� +{,���������5W����j�EכT����AM�J\����J���G
6��&[�gv���k]�p���?�Z�`Q�P��|? �ޜ���>�^��m�%uѿ"ZxY���Ru~%��j��ǃƵ�ӍvnL|F�.�_��
@8�D����C�%}�V��AR���q:a[�!�-�_G�Z&�_�Ai�j�o��{{\����qt��gś�E�S��@���@"h{��9/�ssΰ�MJ�K99.J��q���((��L�K{$:�$��Rcӡ�Ƭ�2t)m����6�\�[���g�cDx��6=Ւg�I��9�����R�ԫ�t��M��l>�Xp��0h*s!�N��L�u��\%�鉻l�N��+
#����QH3�?X@c�/3"?���|�?8!��tŞ���o�B��q�X�t�񑮧�r#歶�Q�h�(��|}�>+v�y<j\y�3�qOm�:ƒR����U����1����V}K�~@x�2(��?�q��Y�yi#�>q�G"O�,��e��w����<j�_n�VfkE����ʖ� ?��To�2?;ڟ�v�0"���]����g�b^����X�-ꥃ�B#��E��+��W.��u����H�
������w�zGF�8��cҵƢ�%Y1;źV�vHА��օNG�X;[r���jJzĻ6�µo�&�B��;������m^�IlHI�Y�?���Z�B�Q}��on�\��2��X22>xs��|cJi�(v��]˕��2=�i8�.!8��P��;��^4�~Z=��&P),a�	��@�c?�{�k�nZ���O #Oo �)�*�&&��aw�}�k�3���OsmJ�5^D'��4Z���0��v��	`�<lt�����o�sH��!�Lڎ��?(-_���3O��ӺJE��&�]�nP%�B^��yw	����^ɦ���p���IT2!�f��	f�����!L�!	H�q,�m��D��Ԡ����c��m0+w;��[s6�J�D���)*�(�� =33$�)�;�xX)}�9 � m�W�{�yT���ga�*]�o�*=+zVt��F�o���]�X���i�	��55�f+�#}E$$����z��O�g���ݛ��r����{D��,�A����u*�a�x��N�g����Ys�B�KG,�u�4�&hs�Sxm���\s<�ݓ�a����aSm�q侢��	 I���Q'c�$(�H
qǖ��ՍE'�<2]Af�γ�5��jZ2Q��g���1�+���U�����C�=�MW|q�ΒcY	��v�h����ؚ�%X�B���L>>�;rS�V4������u�w�&��W� ��+	�o-�7F$�$-��["��bP"1sX���nx4����GڜA|s���_W�i����j�|��U����(�r��n�$�3�?o�k5X�H�F��C��W˔��z�U!�e��C9|����f�b������q\��*������J:9�icH��FC��?���VYw?�������m��,i���C�귶�����`$LG��'�J(�o3�bH�x�꼅1�˥�=d+��N�C�V�9p��I�2�{���,��E��Yq|I5by\�Җ��k9��	�	D�b��UQ���Ne߯'�v����Q$_����j��Y`%�K?/����%e�6�QX<�mw6͈�2��5�j��'��1�x�B3���8𶪀���4��< `��A��w��2�')��72Ob�j��;Z)�<��f	�BA��p�#5]-����D�Q��������I+��2���zk���7́.���Q7�x���7,[�y��Z+��*]��(v��cHb˄�W�_yL>_��0�Y����m�ش^jV�M�x���)�M�M�bnlJ����.ܔ�K4�|��#Μ��ꑝ)t^��q�DH���RH���b���ݭ9�ͼHAk!����8r&t}x�#��ϥ�څ����m§Nw�_;9�t�AB����K�D�rmI�Γ�WǑ��6�>��y�r'�'X�<�f~c�)�$Q����1g�(Yz�e���a�DaZѩWD�P�v�O�|H�Q�Wnh��>|��d���z#��T�Qe��u���`��	�!�[���Nǣ�ȷ����r�x=�E���x����p�$4sK�fG���cE�a�8�t�����&���<�8B��lm�=��h,�`dQ5���m��!�VJo���-�Lȅi}Qu���j����!DN�Ti�M�qpi^4�]@��
E�KW7��hc�[�K