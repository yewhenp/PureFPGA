��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� j^ꘜI��e�cA���t���D���[\�Z6���򐝵&�<�r�
�O{���!�R� �s�W������go<�xĴ�)���5�����X\�H�
@'0��p�?�=��6��B�{L�.����	 ��/�;��=��W��ajQb����Ф�~��M��GP{:��hM��^�}��`^�2T?6'��ȷ�ir:R� !�"��������c2j�F���cٛ�42�#fsq�#��i�D�H���Zy�vA�:88:�q��<$�j���=n =���K����JJ�2���s�%�b��;ߚ��������s����D5k��]@�n&�Ed3�=>�k3L��m�����OĥK��?��Ul?E�cOrZhH}p�I��u�b�?�}�����:����j)�J���h��5�0�(�^{*;�0�n$>8��M�A��
`��}�gҿ�x�[�U��Ւl�n� ?�g�Jo2�0�kpu����A���E&\8
����x�|��r
)v�f|]�� )�^H
�4�<eӓ0v���)/�����v�1E���A4"�6}~,� [m,ॼ�ȗ�C���#�?�O��Z	��:0�RMr�|To��o¬��Q�ի�|d;��*'�w@�B��xކ���#����ʜ���t���¡[��$3���W�ߚO����2N'�H������<���HB��@�%ß����ZG{bN��LfS1LÆ@�\�$do������������+a$� Wɸ����n�ZKh��*1�`�T�=�0��S�C_�t���u<�x�/�?�'�|%�sw���54�K�Y�I��p)�f���yu^�>������fN��|��5 -��R����ܨ�����2�Q��Bm�:Xb}��r��Ep�A���0{�����3�e�cJcT�a���Hx �5��S���$T�O({I:�'̯Uԧ��������7=�!W&���Ľ��m-A�~,������D
V��)q���A<(�P�Eזg|�s���A����^[~�bۄ<�7o���W͔K���D�i�p����j<X�.$����f��|�/i�D�Ep����B�%���ɼ�L�å�*�nTIJ���u0ׇ��Cd7���~]�������������5���ǥn>,��m���7υ� NkXMX5Tb �7��?	��A���)a��Ǿo"y��Q����I�	����S��$�S���y��Ê�a&v:�#.�q/*���H�Duh|�Ƣl9�ﯡ��X�k����y�&KR�Sa>2.�!W���׻��sC����ˎ�hEh����6\]�a9��"^����5�$t �y'��Ā��Y�U��/H5�Wە_Nm.\��j 䄓���i�Z^ |���]�|�4�(/k���R�ڝӜk�5z��`k*��[KU���g��x�h����}���*@�Z��Y�K`I	.�����8��2fG���㳈��R�M[<h��#�!��=��H���c�	����0�����_ۥc�-.���������S��5��Sy�3aS�k� tV*̦��q��2g|�wF{���D��'��x�TW�eB�PXuC#Α��:���{���b��
,��tͨ��	�L�ܻJ\�j5���dyݿ�hݙ���x�v��T6�mL�WI������H���y@��m�������[�Wԝ������s�]p���vW�u�,�̴�q�+R���ח�I�4c�p'�m�؛���o��
�#�����G.;��E���n� k�h�s�w�镡{�+�{)�}�lpR��<����%���hM��2
S�a
��F;������~a���O��V_K����@k�;?#����B�HlTY���P0�x��b�(V�{/8��8�[�!!�QmOUfXx(�ksl���q$�t��^[5�ňķ�f������a����k�*4�<�|���s��׳. �}����I�p���6�_�	O����DI�M�������ȪONǄw���r'*B����r~��C�7��ot�������"Nn>J;���"�Kc�'�D5��2�y��v�$i���zB��a�fb�M���{U4ˌK��(��p˔�ҩ͢�e����c`�n���Bʔ��B�y��s��d��;F�)�� �L?6�
CX���&6hwڕ��6e�u#b{3��7�[63�̃Ǖ�7v��6��n\_(�b��u�V�"$]���׋[����H"���ޤYד8�eE���p	�e�Dٞ6Z��6R����?h�.>v�Y�k@ت�0.�q,+�L�`_�;��*��=} Qz�  � vo� �I�^��5�ø���w��z��J���{�;���͋�'I�P��Pt���~W�pF�[�at�F3#�Y���Z)��ѩ�P ��C��z�5��뒴�Q�� �W�}�F�!)�W���h�p����<����_���Hq~)�XA=�H��U�Ԩ�,�Ҷ��
��rn�����(O�;�C��9o����+C�*�Rk�@��<P��+��಼�ڤ)�0�2��^a�`�*���J��v*��Ai��V'��t�lk�!�JMZ���[/&�@�wҘ�l���K/h�N�v�G�[1|)�J��-���qH�KX�1��T���uY�0�������R"羧�>����p�oѷY����${ܵ����F㍿?G��¸� �;��D���Y��d!�+-��'p͟�<S����_�17Pyk��b�Da��F�S`.��ix��� =���n�=S�i���?�Z���;�m��%�B)���&dO��-�Y�L��U�wA���u��� m���0�,�{��Q�݋�B����rQ	�X�($��	�;z	�edsԂ4J]�B��钃��\� M��[%p���OĪ&�t*��.�����u〉�����]D��:f{W�#~�������!R�v��2�ӎ�^�/x����[Gh�j#��^�n(j��r
�i4=6=�F�ݜo D$�(N�B|!��X�j+~=�!�yؼ���>�֭� �gΦ�XmN�}����JI���8����e�nqC�zm��o��悺�g���C�+I�ޯۯ�eO��qp�t9r�41�X�\�È�[���ti�e(��Ѭ�'~�h#k"Fn��E���~�M�%G���D"2��=�q��c��r3�N������fs�b�j{Ԫ�*m�[?Z
�q�d��������<��<NF8Dơ5X�f���3��͋Qi
D���:aNHy���[��k�f�C{p�6u���g�#="ܯb�7P��g���]21g��DK$���G�� � �:�SYV��2�D�&l�Ƒ�p���:R������6���P�4�u�K����a�S����#��,�<���/�F.ZpL�sO�#MPQ�����w��>�}0[��B��r�u,�����/_G3��f�z�r|�3,Mv���i�b$M��~�!8o�tچ�m����7��5i	A��Yw�2ۏ�§��N� $}C}occ��]�X% �
�jj�>;�ݧ���d�{`J�>���A5E�t�����H�WJ=�������D�;���ԗي
k8S���X>��m��W�=���<ERe#�tFC�F�V-,��^]�}��p��ȗS�mi�D����5a��%�9C����gJ�~��6��(ݒ�Q+�YD�^l�x�D���=�0�C�k9�f<�TfW4�s��gb����~|I�Ϫ���U�I �y��6�����Q�qz"�f8�H���r0w���5WA��!B��ʟu-:w�es�&�wf���@&���\W _��v5���M>0�X��Ͷ�����U1G7�v��Ӷx��0��/U�a�s˝%{An��{��͟����m1.��H�����8�]tN��C,�̘ə)>����ǚ#������U5��ȡS N���c)�Q+<Npd�N��_��x��F���&��*Z�/�J�ʛL; 
p���l�Z���Q�LG�[���Oh���zq���C����h�hS{4�Z�WC��f����F��z ��T�J4���#���W�+\Vf��e�b~�b"�:pn�6�%�Rd�8��Ё�5Ic6&�h�T�8u��B�X��"�%�k�K�?�E*������QǪ���)Fx1��g|֞;�LK�oE\S���{�c2��b�V�}�?OA�lK��n���\v@nTRp�����5e� �N"o��� -[�Q�X��Z�?��j񑚈�m'.g�}+��GiOɯlF0����rfA̭���h�L$�{k4V��N�[��J�%�j���:�Љh\�&_���2�����T�[����<��� �,6w��Ṗ3��%NO���e�aC�)O�ԡ�5�)�����Z�����y$�ߛ��a��|+���*b[L,�Mo�-|?��ᴶ����#1\5<r�̎�>|3&ȣ81V|�3����kPpS�E�Rx"�^A�8V�8���ʠ�?�t��DVI��=$O]��۽^ޙ1�*��u'��.����`g�"BdS��.�+䨍�d���ː!>��׌'B{��n8�����	�����H�VEX�m�_���ƌ6�*��1�[���>�I��븘�o�7��(�H�|�'�;�i�w'��2� F !��o�D�Ǫ��ߴDǇhmS���i����mھ2	�$�B��T���f?c���]kN5�|F]����fi<ޏ��?�R�>�>������?g����\��{�ko�O��vHF��"Q,*��s�t�u��9040���27��ʶ;$����Y���t |AeM�mQ>�5~Z�ClN�cm➦�}>3�O��	nK:��N�~��3I�E�%� ���h/bT-^wJ�/|������T8��O�À9�*D���O>��acy�_�ؠ������T�6���7���3�Y3ed��h�2
�����ZXҡ�]_�6.���{b�!�`����`�&b�4ϾHU:�N���������{j�l�c���MC��H�㾛$D�,��E��� <~�'�A�%5���k��eVv܏���y��� �+�:��5@3~1}��������
�o}|�\�������&�"�����R0q)1�<K���	�N�f$�r�c��!�{k����bp0�N�}�d�4�e�83$-
��jWt���Q�l�)ȝ�$,�G��l�����!���/��ٞ/yf�)�h[g��D�S&5�%�ŰF��Fl���v�@�k��߲a���<�u�g�#{�n��1s��0ݔK�B3r57�����wdU-�-��b��4�(��š�6�ܭv��s�{�7Zu=o9,49�ɷ�D�����{8%����6V��v=е��%Q�Y�*
�,���5����XG�k���1��5N�dYZ�yMcL���k����9�|��o�r4���~{Li�0 %�:H h".�W�х����Tf�[s���F�m�R6¾JH���ifɒ8��^O,�m��&��4U#�5lGǄ*l�BU������SujI8���ƺ;{"�h�x����W�҇?vwGQ��Ԯ��&a�)}���)�P�/��y`�U��;�-���x��%�;�e����i6�C�i�|��~��P�W�UeV	Дtj�]�������|��u�ċ�ȵ�F"��bj�ޙ�G@XF�b�B�MmŌL�DV�`���'ԙţ�N\���n��5*6c�3�?���|oT��p��
`��T8�Ն��[�}�Vig	̫J#��W|Ρ8U�L@�G:�߿����ف}~�5enN�c��Y J������'At�YjQ2=�p���J�����^SU�$MWJ�Ԁ�TJ�W�i�Ot�&-���eQ�z��B�����l�X�x�
��W��:���'� &(K�$�NhT �����:Qss� ��%�4�(y�8���gN�U>�Z��l�2:n�f9��{�ߵ����s��\(�R(]�t�1J����Q�\-k2F�b�7��F$���ޓ�C����d�ϗ��=�7�X�8��0�v��5�H���:}W��Ng�d������c�&()gdi�+�Ú3WS�i��]��y�1W2����"�Hpۢ�_�Z�#{�u>���V��=N�l!�6y>���2}�Y��'A�2���|5&������uVK�򺱽hQ�G�YzA�e9�og*���ݡ�JI���)$_mq�[�4�JQ�ư�6(��C|619����{�&���)3��p�_b��g_�>���n�s�J ~~v������"��Ҏ(j��A���x��It���5��KR�ȩ��&�J1{d�s���?~M7��R�0K{�j���z���sU��Ecj<�Z���ƾ��f�pY)Ȼ�{�@��)�L�v70��RwYn�(ܨ��f�#�0����}���l,!�pt8<&��u/�ז����&�SJ�ʠ�a*�V?r�#0ً�D��S�:1�~��T��"x�LC�O���U~�|
�Æ���L���d�9mC�o��"�>=�W�Aq r0��d��m]��e�yvĔR�<T�n��R���}'�_�JG��:�����BhT��!��;�`�i��s`}\�E�̠�{�-tq�t�f��pA�����A��i�|r��'����r�\�kl$LT��8!J�Y��zX�#�7Z}��;�<℧�����\~�	�0��8L��%���@n�(�ٵ8{��[�N�W����%�>xwC!�TjWw1�=@�� ��7�*~��FN��;�!�'�`�tM��Sd8ǟA�)C2��fڅqLl�f�'����$L+����5擱3���u��&8C�!WrÎQ�:?]g�͊{M�%�9b������u��:�崷Ψ0��xLx��:�5�T��>
:	��J��Լ�i��k���3G��"��G|���|V��QdCH�|SOn}�0+����]v��������<������D�
Y�]/��\�f�زQ�7���e�a�>��=�7����Q1���~3�w��^�I��3�o|��i� �T�C#|t�ξ6�6�o�^��6_x7xi&�e�>"pSl
�AD��y�E��b3�{飕 �����*�ux<t8�v��?yaE�{�����-VeL�D��`�kW�J;/ɾ�K�vbA�ģ��7uϴ<�͢���p�x��{�z��)[xo��~P�~���;A�u�b�h�HE�\tĳ�4�*�XjnD�'�RD���XTQ�5=Q��D��)C\�����o3\~�kFa
�T	+���M�E=��u6P�5�X-
A����[�)��PZC���ӣCTFr�}�nK��+m�)�������a�:{B����8X�Ϋ��.�R#H�ێ7ߖ��d���q@.,�D��G�}��ZB�,��m���L�g,��S�}�����@��Ў4���>ܫ��,-PҸ�&q�q�ƀH� 	3��F�����(�n�D�������;�!)�WC�������C��o ���	�(�zȏ:�h���U�Y ���h�z�#��!��y��hm��g��LH�AI��v����|̈́�o�\����p�VNx�|�c�E\��*�ͫ�P��)(~ԩ��_�T����S�7����-�$��Qh?�q��.�I�'��{^�[���"�,��=Sm�	7����B{�km��_�`0��r��%�4�Ty�K?ۏ��-6���]S���O�� ���H����k����H�A�b4*�=��O��%#%�k�+䂮�T��)����ᇩ��۽��Ƙ	'�Rj���
�������f�H�E{�@N��R�u`�s2tVLT��c��DGA��]_��{�C�D2��2�0�����Y���� S���w9k�Vy ;O�	y�αx�L��,b�~57$pL��g�X���A���mn
��y>�sܵf���6U>�@}zL�=ά�rf V� `���r�-���-�����s(q���JRO[�q�"���L�z}��8"��| J�T��n�&�6��?�Qj9"Jq%*?Y���}�@)��G�VNM`D(��\�I"��$�v�t?`eE�lkjw�"�BWEq�1�h�ϱf}�\�����0˩��Ub�ѯ���v��u�b�f1�W�Ʃ�K�m�o����a*2���� �.&��P�`s�ɇ�o�����e
��^H�"R��r�"_C�v-u�f�>A��X�u��Y_���pK�X��u0���Y�5�'�p����|��B���u�̈,q�j|j-��c-��Ԯv)��7�����K{����[i�r/}���w�Q6\M��F�(6�-ʊm�KW������E:������Xl���hW�,��2+/8tɊ��ʧ�8/Ǿ�E�����N�����e	-M<��2��m����D�
�5����(��L�a�w�s*9Lc�-���g��=��(Ħ��boM�ֳ[��7�f�r%�.l<��C����A7{���9���(����.%�YёP���'H\IS��� �^eRpE�Y�w������ĆD�ݢ4����^�k@��������Y<�G@a���NEiI%�mH4݈�7�$��Xzđy�`�qQ�WC���A)�!_�Y�Mi˗w�[�ƀ,< ����$H'E���g�xnm���e���o{�P���:������3�����H����,�Z�R�]�S�� ;�e��XY��	����(��������k����=D�S�`B�˼�D�!Σj>�χ��º�ݮ��a�F? ~��Ժ���a_u^��$g�w�Xax+�	q�6���x a>?H2rj�Om�|vOas\-W���&����?�E\O^����|v�u��`��t�,'�Rk�hc�w��؞ǜD w(�I�}ěvWz����53¦�xgKa��:��%����-���nYX]Ϊ=��
���5O�?�~�X�J�s4g��g��F&�qR���ƛ�C��X����Ϭ9�h��!_��=��ʤF��J`֛�9L��񹸋j�՗W��5fC�@4�융ߤ���Fc�+0|��+<+�LI�~S2���uz�*3�L�t�Rrmk`I�A�	ס�{�߳�~6;fjq劣�HSwf�Ï@1Hi;�,=�l E(S�V��5�[}p��٭]߽7�>Qoed^O�)�-�-�(p�j�{׍�Z����������Ni޿����V�lzo�� wi�B�q;O���C4 8�jQlʠ�w^����5C����Y^��y�Ɗ$�4���m�Z\�m�i�nu[6�B�n",�(�#j3h��9`��xAe���eíU��Gj�������+��/�0��>��#dJH�^���J+�p�W%32�/�jL��B]��:�6��R0�=p
2��>�
�mqq������c�(��Aqc4�G&5s�b[ø��$Y��$�(�cJȭۓc4��5j��~=���*����z�7b(�D�p$�k��t,ƪZ\uir̯�oGVdJ8S��qg���%N��}��o!pI�Y%{)8�(�y���3u7����H�y�/~݄Sz��b>�F�٤[bzdű�]+C�$v�,�B�F���p񱭯�>�C?uec���Q����7�9k`f�P�c�MtV"V[�W�sPkw�Y���~y�"������H��ݎ:G�5!}��zD��7 �(w��Fu2�%�������K>���4i�en�X)<�H28��]]2f߿��[9_��7ps���S��;�6A�['e���oI��gę�A *�<�%�|��t���P�,���R�4�iS�9��>��8_)�$]� �Э�� Ǽ������B�'��g��D�����+j��Y���F<U�GM�{�D��-�I6�����P̮���Sb�6��jgit����ǝMUjjT#h�I{H�>����o�zB���t��A���� O������6���G��\��4�f���8o��PJ���}T;?=ʩo8�I�Q/��R"�̄�Kl�pʯֵ�g�>AG����a6z6�cɩ��(�{�*[��\�)�;^?�]�}�a�qWs�����8��.n@���N~���(�Bõ(�D̀�����J�b��Fv�Adi�����۞���W��hj��&��|������l�@�kA<��D I3GDkJ��WV�a�#��ep��o*�Ѡ�{�=9�}��u�U�F���$�~��>R�VFl����������)�$.���$��	�^Co���L���Z�<*D!O[� ����r��'غ����r0��� �����n�[F
Iz��#�L?�MŲX��$~ʑ�r�%Sw�$�8�P��w����u{�#c�a�5Ң��Bј*;+�u;@�( ���0�W���������6|�a?ꐌ�Sժ�C���6C=3�唩�J-)�g�����Z/��m��=ri��O#�?�t�^�bQ4[��qv�~���lgg� �I	����M�I'˓ӓ�5�s j�^(NO�e|���׎^����4�F�&J�m��|��#m5��#[+Z��N�M$n73����Q�t;�I�7 w�S���(We���[�b&N�؝�Mq*�m���.8��
�<d⒦-�=^�}9�����z��ʚ��.IHU�����?�r���e6@�� ����\�����to�*s~�<:��Ǔ$���w�';�ldK��&��n.���W�"S���0*d��r�arz"��]z}�<�3P{����itm݀��r�o@Y��6i��ki٤��`�i��i��-�%��8'I>Z+lx�F2��TK9**��Cuc�ڥ"S���,�G>ʖ�i���N_+}������EV�bm���9rJ�pج/�e"���[�4�4�b'K�ϖrb�&�������%�bfh�[���w�R�����"4XߕH��k��-w|��eh�)=�����n�[Yd��,��e}��t�A����x�<��x��[ݷ�!5$V[7bE�X�'���j�u�t����^n�ل��" �:��iU<���׬?��K�l�:Ϊ�B�k��EtK �{�|a��VT��<����*�5.�%�V�3���o��z
*}�6�=���g�ǒ�ˁ�˂K"����I���`�:�$�N��^�:½a&��ň���PΟ�������L��I�qx���Z�[#	h\���ǔ��|߫b�a"�����y�F�榼�9m� ��߈�"��Z����� �	t����z{V�����)�H椐@W�w~ʜ�g��!�;�g�c�AWk���M�%	�p��'�C������g����M�����1�%(��d������1�y�!�C�������6�w��X�rm��s�4��Ҝ�����RѢ2�֜X�Rh���c��u`�W2�hg9So�Y[��C�}�5����pSi��L��$G�R�������_��v_��I���Ѿ W��C���_�sO���q��Am��G��q��<��P��4B��K�I���4!���k\f�����a��fQ�a�3�����C��G^��!��o��6Rx�7�� bq�DSé}i�W�-���Z� &C���:ǝ��D����C��`1��j�R�dd��7��b	�&��1+jm�`=�?M�.�\���L_7l���9<��1~��`����B2��,o�ص��	W!]��.=���F����Z�Z��E���=��;Nr��t.��N�+��e���1�{P��)=���{x��|t-���*���'��;*6E���kH~�z�w��^�!#�`0e��Lj�
�!�5ה~tz���.�iò�~͂�K>�%��4�y�`�*#'����B�3Ȗ�gz�x�8?�e�R�sD�U�flp"'����Y�ş{�r����y�ȗ����ڣa�K���4����5]����%�6Ce5�w�;�z"�l 0IՑxeU�x,�'(�φIӒ49��i<IG�*��\�s_g��T�k�kOG�(�<-��/���i�cVb���j���`߮?T�S0 ̑��ݕ��̻�xF���JVq�0s��F�?�g�C Y�d�M�c�nkt#�4r{E��Z�(���?�#c���1�P��1�)َ����䓯���Q��^uIJ���\�h^�"�v�SMG�����g�L}q���Yqxo1i���9ۊ!M6�kqC�Ֆ4B<g�7���Ő�?��d�$����1�3s<O+��f��3�tFس8WeI���/��-�Ҡ����2�]�w�J���)D�"���T3x3�x�d�r�J݃s����>w�f����K'lɾ�YNp��Jދ������̊$��� S9<����!�����8���C�Z_x����GeE����C�,[��7b�Q���4tvz,�v~�^��	;��"gu�E�V8�(r�5��n�W�2u�v�](�n�YZ��Tby�a��L)���F�i�q����ey^�|�Qa����{*>E/j��`b�zI	+&�	�q���D�*�����(�u�2��R�znl��\�oJ���2���V�n7��R�uA-�Cv�[��g�y�V,:�aHy:�x`�*p���\L��\o����+#���야]��;��o^��ɹ[D�~�,]��E���e4U>�a;E�ֹQ��r�曂*!�9y\�푭�
a���p�som)����^Gl���/���5�nm7�mI��ڋ�@$I��M�΂(]di�J:X�YFE�=����c &���h�M�G�%�_X�8���R�_�n��:D�!�7�.G�˶wq#���w�/8��UҞ�(¡_��dޒ��̙��do� �_	������Z=V���y8�x�⪝&���4�$����2��~����5D�K)���C ;S�L����[�z�P�4��+�|��H�G�@�n$���BYk�ɑl���2�8	99��]c:�]�3:�gt��m�E�AP���$�6�Hڳ����W�dQ��VK���L�J�����3�M���VO�q;�gԊ��q�u�Q�J~a���♳�_�zm�'�vNa����>}N;@L{dY��B��ϋ�q����(�m�eX�6������
�Z˘/r	ˣ�)����
eF��S,Nm�.�*��4�^�J �|�5�G�u��K��Ӧɢ	0����bƕ}/x�0#t/I�Y?\���oA8}'o�9�ԝ'��.]�����A��= �4�Uu�y݂s&����E��ȋV��%�"���j6:%Z�B7H}�e����lU`B���t��~���2��ү�t���|æޖE]�q�[TP�T���43���W`{�+�&�0�n�S2(	�V剚��q�
Ok=�͗ɰ�s�N��/�k_Vu	���HPzӱ1���ɘ��>��ߝh2a����� [��|�E4���krH��<񴀽���N�~ט�Յ[�x��>���I����]s�%à֢�>���[�w�T�8�A��xzRe�R� ܉CLH~�e*�&L��s=u��r
�J.�:�n�R��zC�On^�Zzp�9.�E��xsì1��`(5���_
����k��K�i�uM�(�bq��BPS�f��-қ�_k�#�������[gQ�gζǎ=����S�R���x�X���fb�}�mJ[n�=�V�%�ADLʁǤcČ���@oX�����}F�̗>�t;j��w�z3K�^-8k�K#c�t��=H�MiD3���K�`э��PՁ'x�-$��%���+��4��J�P��t���@�n��j�Xo�N�*C���c�ˋ���F<	X}�1ɂzR
�[�hѰ�%J�eK�^̓���Q��� �CEbq)�:����o~Y&��MSڢF��Vb�����},W1%�i\A1����#�
�~K�k���g���@�9��
ɕ<ԥ����od귆�_�����\B�S�4����J�1�_��x)�D����3��"ޝY.�����4w��T�ǩ���H})�f����������Z*i��5
#�/NX��H6n=e1��΂�w�u�����	~��0(�aH�%���g�<�g!4�:_��%0�J�(��C}��+��1� �r����g��39q:j��)��Z&�#7A���o�&x��{�+�R%� �M�:͈(��f�J��n��Q��Q�b�=��/�a�蒖K�s�|�>�GH��	�o��)��m.4_��WЗ^��A�1Y&���Jt�#�(��vw���� }�A�����At�8��եF��%�����J� ?�*d#=Yv�¼^Z��L�n��O�@U��@}�(�`���7;��&I�B�v��R�Z���e��/i�m*T'��5P\:�eR�qf~��:��N& 4O���j�M�j�#�e ��v�����y!n`��҇�a��:�f;LW�}��,�������|�>�J�w� mCFUZ8T1X�W�B���/�����Z��s��x~Y<��lt�<�d:I	�8�_������,��d�E�������D���Z��f�x�,w:�dt
���ΞRF)_{���,�ME���*���|H���� ��b�l-�a���d܎�;��L�¸e�La5] �}Z��(Z>�z���=ΘZk�c���A�Ǡ|{�1Z�Kc��,ϯ�!�I k%1��q�`��֜=Njd������=A��;�.��מ<Y�C�T=-h��3R��5M)�B<�R����.�0}��ܙ�����c����O>����C��XN�0ӥ��;ʹsJ�E�N�2�?�C�	T�)P�Z��9�����'�e+���<�Kf`���7����(���R�v,����(/����D�����?Z$bE\�t�����;ҳ�a��6@���>O�
d~s�
�h;X����lVg��Mz��$L���uty�}��8���A��>�A�{z,p�{U��E��&�1���7�8�jIZK����Ƿ.sO�Meq���N�E����$�Rq�Vk���/�}�v�\^\���~��+ 7�,����J��K�n��(�
�3��f�/EA' ���R�ٲe��o�"��l5b\�~)uwI:h'11HB���8c1_^��p`�eCㄹW�v���0��q>]d� ���P���k�%c�97�]�cw.�]��v��b�-�Kv�̂�c:�>�/N`H*�n�M��5[�n�{Y�f�����pnw#J��`��Ó��86!=�V`T�k��W��	b��;�z��n`����0sNX\$���,޵b���>�G��q�ҳ�}��>���۷E7�kƌ��8���4�C���ݼ݂i��o�W��a_-XD���3��ąl�"�-��MrjA��+��ᚤ��s��`����Gܚ��?� ���g�4���9�TIê�u�d#d�-�rWt]����h�r����;��ф����UQ˨�1U�J��B�)��I�^}���3��B:���{�iE8���������}�ZI���ƙeUS��.#����)��ٳfa 7���z���R��W�ޖ*�S�00�!	�4<�w5����H�>&V ��HEq�=���;�Ҵ�&y�;F�zgF�F��8@�j������r��wq�������
	��� �=�&�H�R�Dl��+-L�����ǚ��@BMQC�q�kUKz���O�S�k�� ��)x:~��}��R(N5�ʏUI]��w�x�C��� |a5�g��\s�� �89	�J� �
V��uE1+��*��|�d���P.�ܑ?�}\P�:��E��n�P�Zz���T=�Ղ��#r�I.�Tn��j�t������j��3�t����N9��`�i�=c¸7ǃz쎢�Ɋ�"�y]���F�3#�2�z�P�qB��}��6NZ�W'1�8
�|'��lL�����L\�R�/(O��f���!�����!N�%�L����߈s�`�$- ���~���>A��ē�&C8G���v������rڼ��7e1�����#̨� S�'q��<~M��[��6�:3�s�Q�Z�w]*�^B\<�
+ÌV,|��p���i��RM���@�����VG�I���!�?-r�'?��/&��	�) -� U�G}���|A9	��6����-
+�
�5�s��޻�oo2T`�1�prJ�y�W����#�0֠��GU[����ٮiصy�Q���'��j�|�	l6���$�;u���I>S&&�d!���@�P��3Ӝ*r[%�rl�����is�R�æ�BAN6��:ɇ	���l'z�(#{����LH����7C�>��3>�Ͷ��yaa��hs�R�N��B�����\���.�L� �G�N$�C��whw<�~d�ݷ�ffZY1R�۳Ho��S�Or���Z�%�z�j���0�r�?t�3�|�?�.p���!��z~_Y�բ��A��k��/�V,���0�j��v�m��ckC�ն��Դ�&�O��hT���:�=1Vx�^�.��OӉ�_e!�aM��7atR��O~�p�����#��'�_�_No蓲�� tr��<WZ^�;FQ3[�?3���Q$3s

��Ҋ�j��у������+�N���f�㹖��|c����i�*N���=�~]� 
hR.g{�Q�JT&�+R$�u8�p��
�&踛1)�2��!Q�K?��u ��4T��hu>���
y�xa�
��	�X�?2�N��`�Q��bn����\��3�D���6�c�c>@�@0�$��-$J�B��/`�Z>X_#���0��kd�����!����.���)'L��:y�J\�]�v�|
*������%\9�.s�E%a���s����㝚�F�{P�]=CS�s=�h��a�;)E���%5k�7������h��<��އ�yFg���zYQ���� �΃u��:&���7��}�R�2N�H�����c�{,���mۙ�T�rVy��\5b���7�n/r��T|��pGw*��� �7m㧔M>����D�Z�<�= Ƚ��M� ��0X����J�Z$�框��8�_�l������bp,ц���=E�!��ḿ�Z�nY��a翝D؃�R\'�j�-^
��1��w�<��Hg�u�6����8��SO��v�l�]]8^t�9�h�f�C��Gddc3�� 2�4�W��m����R��i��Xf-�y�Kڝ�ۚ��-;�զ,��Rǥ�(�ݘqy��˖�%.���(w&ҡ��v��<(�S�u1+�Vg�df^��
ec�Q#Kнb��ꍆ[��`�
�E������0�0��Hƙ���3���8��T��s_����<�؏`���i�X`�ň�b�(�脈9]UƋ<Fʂh*v7H���j�,���q�jk/�+�oȘ�"wB{J�9?���w�oP"���%k��9�Q�5�q[p����&Xj�п{����l�4 ����k�eH��A J��������?�zڏ���+���� fK�_i[c����\T�fRX6���Ѽ��M�zBnf\�@,�~����]�1��u�4���C�	�'�k�l���XHd���]`�|w��i��o]4f��q=� 
�u�P����5l���@�P(�R���6Ѹ%����NE~�W�/�h�4�y,uD��Z�z��v}5���ݲ�x����S.8Z&<�>�I�v���e�`�@��_إR>m�96�F{�	�_���?���(��*oՁ\��~�e^,W~�ذ>�z{}5j׷��/F��C��ٞqfx5��~�Q�y`�0�3sI��	��4�]=��s��Y0�I�N��I��w�������,%�UL4��q��6����1�/06��\��@��Ou�[���ر��ڨ�p呬�^A�Ӓ_a�W.�4��2cM������!�&��
��o>��(1�W�F�n'�1�n2�l0coI�I��o� �I�&N�`�b��`IA�敆���Չ1���(g5�.g݅+���.�	P��T���ۥ)�}0ls���B̌����D�>��]|�}��<�.��+���R���R���������ٙ���>�1ʚ4W���+��M�.�KMW
��9kў&'%�RwQ]9�30�L` {vsF��&tN�-�V=9$+���E��Q
A2w��˒���iQz���y�����F�!�5&�������p
���g��>ɴ]t�F�<��]�)���W�ܤ��uJ�V��NC):ٲ��/���"}��t���)��$�9�`vE�R����n������E��b��c��چ����<(pRx�nb#/�?����.I��W�E��_�3vc�np�����ԍ�VֆmF{:�4
�PNbj>��E)�쑗I�����V��M���C�^2L�gY�8c���;�<N\A�\=���Ó�V���pm#�/9����jT�:''�"	��IȡP�ImG�A����K����Eu��"��Ԍs�+�!�a?��h;(:ޜH��}�]�]�c�Q�4�.bT�~+�z;B,�UI�"P�k����9A�_�����]�F��=��*���N�1��;t����j,a�^�p�k��Pu���&��W*5c�!�GeX!Ғ�K,)0-ze�_��8Z�f'+\��+��X���Tey�у�'���{��%(f�����8��:+~�`\s-7_.VX�'��u���J�+�O�o�l�KP!g�$���M�A�n|/�6ӭ�����~��y�Ô��	E��=Ǩ�-/`)�g�lUm�Up��'|�^�D��s�l�����Di+��>��I<H:�,�.i�W�&�G8	���r�^rwU���:"Ȋy����Iv!�wɒ����.�O~���q&��������-�wA��@y�����2|����ơG@-�Ä�p�+���N���D�Yp�A��6K�&ɘ��¨�|�������%�[���%�yWv��ɛ�V����ѲIЍ�������#��>��v�ì&�^�!��F�dw7Zn��܊x׿�DS�b��,�g�z�a���@a��������\hQ5�q�͡qC
NVv���ھP �V�߮ݯ���kR�����*�x,�;As.�-��)�v��D
Vz랑���<~�Qj&p^�4�X�����E�J��߲`�t��"-�7{i-q�e�QQ��
]���|��F�������Zm��룷�B�y�up�KGh�3R����C�G�j�x������*]��䚺>O������T���#�S:P�?�ȩń|�cg�*�k��y,q�h�ٗp�"�[8�q�6�:(�l�0I��75��I:di�@�=?b��n�� ����+H��K)z]�lw���&��|ln�H���K���X}�nz��%�)�7��f��2$Q���fs,��.Lt0��M ��!�������U*NWqpHx��|�f��@��/_יt�,%w�2k���4<*�l�{4Of�P���"ȗ�-�eYY�_��5���Ll��/��u�9\�	�sF��%���3S`}��h��pPtÛ�����	��K���7������R�cz�I��A�Ani�Z��?�%�ѩ��������9b5�0�fq����T�	�u�~K�$��Wx+=��^J��7�g^�G��d��8�Q��b��U<1w���v��v5�����o��b���8E�č���9�+��߉�@���Ƕ&cI+��n*��E�G2�'X}�U��Wl�k
X�y�y��5_2�*�z)�4m��6�kO�����
<��b��r��ԁv	���XO��ꛔH���젆ݨ��@�v�<���z����`��{�����Og Ȉ��I|Y��?
�9��Sq�W���D\���.-�{�ӞKuK5�n�	V/���Ñr��
ʸW�m�
n=���G(����f\x~#���:�搲��zݞ�UPD -�O�X��{������ �]��U�>f�ϧk��Y��y!�B�hUJ�yq��I�����M�,�urRR�ݵ�̸ʁ�	<*����Pܞ���Q�
yL|�p�t�:v�<٪7T"��r�k?�$�k�	����c�R��nT���Y�t��FXFZ/N���[b
�`�*��&���+(�\�oThL V��K膤-#�|�p����
����RL��l@R⭈��(oo��f���q'�3S*M���7��;ݡ&�_�n �-9��xi�ǈˀ���Wz�U55j7a�}�	R��P�x��3i� ��r{ZZ~a }������d�/��s�G�ԚI1��1��z���a��	>&gz
u��U�Z��V�v��
�I���*�z��k���N{�|/�=�^����n�P<P�;����L#����W����Ҁ]�잕%Y�DBB�/k(��\�d�dC�޹I�� �K�?�Y���	�(��l'ER�rH�*�r0$"{�,c5~�iJ�F�j059�(��d�m��\_-��\\���Oc.���#�+�uؿ��U�|��1-�~v�UG_��̸�5k5٘�w���΋�����7H SY�j�b��U��N�(�]���8 p�n���P]7
<���\��[��8ʀ%�v�%�1]�j��������c���e^t	�����v�L��튟�ד�M�P6�#L��Tݲ�5��*ڏ�0�4�>oa�%����U&��[�5�<��� �z!0�<�R4����ہ��s�, �q汴g\C�rb�>�lEPW��l(kϔ�Q�v2�l���{�m�M(��Ƈ�,����h"�QdJ����^՚��4R��W?P�k�f�hl\�Km�D�-��9�?Xk�M�.�ty�|��$CJ)���ʰ%�qWӾ.,�,�N�,�귚A���9Yb�̢5e8�T�T�$�T�J;���T��&?�t�,~�O����^VD99�Sf����V���2�Mў1��Ѐ�=����ȊyZ�k�L�ޖ����X���� �2.ҟC{&����@r��}���$�t����$�UJ����4ˬ��2��0�~�0�hQZīwM��qK��VBJ<��e3����3_�IG�6����"_S
V:X�����<\�����o�n�T,i7zdX�������=��j��t�8̶H8�z`�a�����{�M2��o{�����sھ�����y���ú���������l^�3gA�8�I��洎�zd��oĘm�خ`~�W�H� d�mO�>'�} �_痿��_!(~�!6�i��,���<o�s;"l�N��Έ�=ɇ���5I�϶8��s`�(2�`[��K	�x�������_�cgQ����9���"���}��U�y۷ɮ �4�e)��7�vG���|9�&���8��MS����Ї�M�p4r�>��nd��A�s˝��`ٷ�����<���3C;"��Y#Q]� �yS������i��ϩj�[�Y�;$�DlVv���_U����~C�ɇ�T��H���C7U�U@+l&tq�mO�9��\��4WI��D��d,b�u�⫧W 55׷W����BZ�G���Ѭgp:4��EbeTG7ʜ��t���<�I�upm�0�KŇ�����ŷ�cZ^`a�L�6N��?�n�M��Vە���u��7�K3�?�O?w����~q�y|ii��)	Wٍ�V\Y��U<��լh�P��Y`�!�E����F))%E%u\��Xz����� JŖڥH��4Ǖ�3���Y��T����$�̂QdN�PG>������
N<e�^�!6��Ws����u�F_�764�Ol�9�xڇ�غ{c�L��kY�ś���ɵ�x�_�]�1 +���+yc��rFx�/���W�����?[�'���zeoCJM�2�k,5C���!�/�z=U�#kgJ���E�����{]gB�"<�(���Z� �,�uj|���޲�s!t�F�ZV��O]ܢ�z@�?x���J@�N,�8]v��gNf��0 Gؕ�*Gw~���!�n.bI~Hn��E�(���_�\y�b�b3���8�n��^�߮�?S�}�S"�l�ɗ���X��J=�&���y�NG(lݪӈ/ꅆ\�������R6��TF�g];L���&l>؈�Z
Q��3K�HP̙�ȣ�0�}I�V7>eC��Q���G��`X��{v�Q���콡Ģrm
�������sț�$���ۦ)�>	0ZٓH���P}��=�;޻**�CӦxφB�_�����[���e�OP�<4M��hj��X˲!�r[;M�4T�&���N�|J���v�J�J���~j�fM��D��,��D-]0,��<��<R��1Q�d�wv�4�U?��z��H��o(�H�c\�h�2k����jCj���eǫ���_mC�Kj�_f�?�n�<#��hU	��/��k�|��v��n�s���\��}NKSN��{(A�$�	�j�eO�l����*u�a��F;l�3�����߻V$��39E�N�c	�>QJBLG��b0�ҭ�j���~�W���,��w���ލ4��$(��(|[��H0�ڀq�q$�=oax?sNkK>~�����	a�Yr��9��Y��F%�=�Q��Y_u����Ί�I9̮e>��ߞ����Y��e;*�z���?���me[*(s��W>B�'��2R�ePW�dT9\9g<�f�=�����O �8�>`�'���R
̧~�п�n.�ױK}����HPv�ƀ�M ��&�M��jvq�����9[����j������/��k��V�r�96m�H�� k�c�+:�������"@�VC*/�n�c%Nfyg �9����j���g!�o��ehY�6��%m��x�xв��C��,�~�Dz#�R8��$"�c���.��bl��ΞX���jr@�Y+�?���N�K�o	����KQy�����9u&�p5��L� #�*��-p\�C�^�����U+qtO+m=�)�L7d9^�t��L"e��x!b�%6�bP|��ک,P��K_^���(���uv��r�I*caK#mƢܼ%�S�ܐ��%�x<ILλ��D��]6�����/jG�@%����?.(4As��Ԓ]j	�*��񊪧C��ue)g��b����m�G��?4��a��+��h^�ߟw:���T��ш����z��*�2��9��l�;������ַ��?K�\����~Kp��R�	<�b�j5}&�{w���c�$c8']<  �S�E�F85��blqdW[^�HL=��!S��m�r�J�8�UΟnM�mٴ@�L@uzB��Z8�_g�� �mU7���1��j��/9��yZQ�`=i"�&I�d�P�]�O4${�X��8�4ݓ����ߖyz-�Qm�fzA
&E5I9�6�P�&2{i�����!/X����<mI�O�;;JE,O���Z`�>�@
H�O�֍M�����3�I�yM��D8�'Y��e��!���~�?���.(���^�z�K�\��C9�4$3y??�jtɠ �[��Ӥ�EX�I��\�T��:��u�"t&,X��À!�QP�p������E��O�M��	�?���Ƅ��+�6��"fp���|\����L�!�0s*�����v/�f���YW�H~��A��i�N>݋(��lD�aU�|�˷x;���|�L���H��m��&�N��<ʧkL��'/��k����� ��`�-nx���7��+�����[೗�,bB�m-h)�%����p��~ ���K%����s��V;���a�����+R�Dct"=ɀW�z�=P<dW�=H�k��0zB�o�f^ �<��C��B���&�ԣ�A���5�����J����
�2�XH����l&~w���*P��s�b:� M��"޵��?C�T��c����H���A}
�O~��q�c2:�F��q�e���\�ļ������2$ʖ��g�h��&O*\�v��@'_�q2��+����-�+����6���B�1M�nk)��yo �X0�0j+NE�.`��	�Y��7�v:)���,#g�uD/���غ��W����d�Q���|�k��D�Mq��,�x3Y���D+�����J��ۅwLH��~ʆ��K~\��x�s`��ə��l��f__j8_�	rA��x#Ȣ�q	�q�7����h�9�֣=С��-CX߹Q	�B=Q@w�-����p��JH��L��^˕�N��?���o#j
��l��e׮��kby����cdVu8\��r�>��r��,�����r�I��� ���?��� -8
��՝�r��"�����h�D�����NucXHW���B�=e٠3�P�DM�&�K�P�q0Hqɣ�^HB�G�{�z��-�e˄ˏj�� �+`�}�Μ�d�w��5Z���̀�:��*�����hv�F[��H9���s�kڔՊgQ4�~��v��蔼�?�Q}��ǣ^��.L (���9�=ڮ�Z��*�!*Ȇ97�z �������lVM�*�1E|[�!��*p��T�&�K�ZR,�p��1�Z����'!��R��#"���)�\���P���EP7�)�����9�H�X����+E�ؕk��\�o���BT�6L"5�OK2�Rd��gA��!۳a/�}x	ޏ�����-/�Cߕr�@iI�U�����BD�b�<�O���^���C���K�Q����?BnU1��p���,o�ȟƅA ��yE����Ae;N�@��Ѧʬq߁����G��J@neEG.�3�{��b*�_�Uau���la��q��x^p�|�KM1�{�a����=�KE��ՠ���ңT5D��e�D��s+[i���&�PEa$�î����9#����|#G*03x�����Y����ܰ>:
���l�D�f���ֺ��x��J*}��#�9[�]��M��:�\��B��?-�#k*/�~Wi)���`sP@�û����kl�6��e�g�]~��If�	��� 
V��d�Bh�N?ϭ<ي�\v �p�k+���(�A}�*�� 9
V#|'MY���'���;3��J�����{&*ۊ�ا ufY9�k�|��ɇ����V庅���X`��D��P�u�Z�-xAD�ȾP=�}�c[|� �t�M��K�0Lg�����c�.K����Ĕ̆��,��'���}��O���(l����r)]k�5��;�\�s�k�+��?9n�