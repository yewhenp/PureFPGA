��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m��k?��V��6��"�"?
���Uڨ�9���52��kD�( )wNފ<vs~~NAuU�k�,�&�Y1Oxp}L]h����b������8�Į���9��r
�+��:�x���8�҄������^����&���e���v�]Cؠ���2]�-m��~i�+�7T��lZ�ZeS��A��Q�����EpCV�7KI��X�4�3_=�Z:'��ͮ�aP���C$��ˡM�vP�%c����k�xa�<1��>-i_?ϩ��v��Wj_���n"���@�OSV���t�k��v9	���>������gd0���WE��ʗ�9�c4����=&�F��� #?���#��� ?�V���l��}��񂺏a�^��jP�f��\��-�qà��}��>j��+(&OT�Irĉ�������D�1�Q�Ig�6b$�n'">���3IaΕD9�� i�ttz���]��C�И�����ЇK�G�j}8M�Y?匛�;�7�4�gP�-V#u���|����kN=��$h��\ݖ�u�Ay7h��zf���$�9Fw���Wy�*�y(	O@d�$G]+��-�����4�����ΗV�ú�d���'�36>���R�iu��XE�� !�C�W�}4 Y`eoZ��a	b��J���I(��)T��V�\ȗ`������{�D��`p�f"�<�zP�%����Ƅ���œ�4��/Yf
)�޸�0�YY�x�{
.ÿ����$몇���D�P��eA6���s�]�I�%+����� {S!�;D�2��Q�S�Ot��5W�Q�W'����Z�<ܱ9@�@� ����f� ?���[�4�Z9'
����U�]ՊϤB��c�z�;P�1�l���������g�?�-h~kkh��'@8qs�2��ګ��k���4,k���z���gw8�|U���(ʤ���>n��t<"B~��#���\ȗLa�-uD���a�?��sKAM��si5D��j62����sFq�
tE�h��捔:��	]�`�[O��kOw�����N�ڽ���Ey��W��w���I���_(C:�v��y�z���ᵍ"�u�N�}�
0 �0-HY��!� ��$�4¶����[���o�ɬ=6Y3��7��K<?qӟ&�V��VLt��(%��k��
ti�(Fv��C@�ej��x��j~����se���R�m*�D햷�ʽ1Y]p���M��b �X��*6�u޿'R�|o��<�J��i��L�>E׍��V�·����I_6���/fYR��*��5◹�o�ژ�!,��{|>�f&�/�D�;���R	5���>E�C��� �0�p[�{���]̽Θ.��O�>��+x��H񺧗����ןK4�
�����X�_j���d6��6���u$����������T:����&������Ւ�g:���*� ��-i2���d.A�Ze>���JK?��Z�~*�	"�o	�͸I�;����A@mG���ҩ��5�/ح��VP�����r�	��Eٱ�-.>vj�����:�e-�5�������3�~n�)��b7{�֥���cL���h�mn��-k�7�fj��+~4���
N��+"����F(?�3�2�A;o����	R�<����>L2ޅ;�����l�J���^׷�v�A1�i�0YG�y�{������^y�ζf��&����Ljn���E��t�
[�ܶ�I �?i%����=*:<B�oǺ��[�2��O[~��ؓ�����[��'�ֵ󉃕����XTeH�ԇ�\�U�5 W;T79	�mBa�p�B�I�}SD�t.LM��{� �P.��x���h:�o;[N�(���*ƲV�L��ǖM1ގZ�0Qƶ��\vY�V) ���.�����5̘?���Ե:����_y�H��j+hT�WIɩbޭd��Ľ��A����G#����G�� �JX�C<j��!��{}Ou~��	l����n�Ɏ�� ��w�����b����X��>���������h�yA<;�8���K���R��3���3�Ĕ�!�������	�XR�s<�Y%�)s���/�f�$=z���tINp9�d���}�[U�mO��2�01���#�R�c���:��n~�4��߄�L�:�����Qv�Ky*m��M�Wf��j;�
��c9v������B�Ш�����6 �� ��,�����8`ǿ��'�}y�^��t��z``��W������a��(	����*/�_6�K �+y�pP��B˳:j���|ڛ��o��?����]���V_�{�b$Y1�қT*�UG�K�����[9�!��x=['P�Q��ƤC�oE�>�+)�(5 �L�"���1NE�V����MP���b��iAc�j�����5�u�:n3�1���� y.��E�,+oⲛ�R�B��i(���)m܃�H'���`�D'd���G'c9����b�0�\�Q �)�Npq��?o�`x-�K��B?(�N����۰a�&��ҿ�? �ق�^�T��9��GlFfʾFb����!���M	3����䜗]ѡ�f7N2y��Ÿ�����v(��E��dޫp�Wͫ���q�3�U?�]�$@�U��EW�Q����"7�/|�������'3�U��!���EU��:�s_NmC"��x�����!��|�x������?"�=o��x6��HhS���,��-�>?١�'�<��!#U�y�m�xf,�n	��ƴ�yn��q�#3������mf4b�Yq�`R��Vs1(�o�28�¿�=)��4V{D5�t�wF��Ec_���ΫuB`�+g<��,s�ե���䒄gr!!�`�S{�>#�^��7ȡO���_熛d�yp����cϓK��6X
}���R/�󏑜b�?=T)�}��T��n��=M��38��>�Q�����.�`�̂�����rV�D]�}���*ږ�^�0{��SYu4ieQP���'[��ȄRP^��Z0I�.b���]ǰԐ/��K1a���e�R=��F�eT{�O����O��4o�R��t|��W����d�ֽ��ʩQ4#���ٛV!��<a|zZ��6"松f�ԩN"��\dP)ӏ�Y�Ǌ�A�JJA�ɺEf��7����od��{��i���4d��_))LN><o�s7D[��wpĶ�M�����e"�e���1�V.Q-/���)lb6�b�ע���:��6�v5�F��6شw�C�x����#��;[� ����J���]�u�Vǥ[䃩'A��
��3�P����$���	��v"�ᴒs�MO)�yd�o���H��]�֣������3���F���/��MȔ���Ap��g�О��P���� ���QzccCE��|Z�X�<�WTJ�<6�G����T>�^�Ԉ7%-�����#�ao	+4Xc�!��>��$9��Sy�HL�Sa�������8�������(�;�B�����J�7n�q��U���)�l��$�L��6���/�Ĳ���aC�NWb��5˴��v�~��d�d�ˈ����#�湇� {��3<+�ŞG=U��l�Ϭ|�Р��N�|z���J�AA�:73��&,�����g`D�`�7*�%�t,��� =Q6��H�� y��V�����e� u��ǭ]\Ft]�Ē�$�3�E���뇹^�1��(g=��cRKUA��1H� ˘&sM�q�S/�q'��f�~�-��;q��zbP�W���|z'������d[`�\�;�k6�W�f�ľ��a����+�����sT�
^D���c�y�������+!���\*a�0���mА/���]�H��MKO���܋��@����_U��|�М��JFp�Vm��jn� �7w�,�7�L9�2S�� �"'�%�kC)tv\f�rh��]���'b�ϔ�Jm���`�IrJ�{���R���(�I��9�S]+M+��3����@�b�	C �S*#ƍ�Ꜳ�X*��D�a�,�� VX�#�7�W��<.��s9�9�lՔrͩ=�������+>�=V��-���
�h�e�f�ބ�}��>@.h�a7��K4qM��k��S7���#S�w���.��M��z��uo��,U�*�m�n@��=7Έ
c���D~�߇��,�ɸ�Ԓ���,kx+
�%�k���L�����|��ܫM��P\�Շ�ZH^�M�c�m�}:��9V扮�Nt��J��W��-��:+f- �y��]EB���M���Q����[s���@��d��NIm��>�$�":�Js5�`鵺B|q~��� �AO�~>�Q��"AP�=��W��r��P��Gp��Zmrx����M��!��~�G�����(�v�sVך��/P�,;r�Uʐ�Yw~���[��N}Υ'��d��qU�RR���=ϙ���h
Y�BGɍ�Huʯ��Z�Ɍ���o�)	�wVh,'�"I��/e��v�5�}�B2�������&�N�������{�y��/�Lg!/ۺ�٧������*�Լ ���9�0i��D����Kj[�4�o ��@��8߁C涍�1�d.1wM1P�(?�J��y�B	�y��m����pT�$>��-%a�(�-��B�xS9lg����n2| ���5��[� S}� �ȝ(�K����P��p��Ui�4-�d�_�"�l_�dy@	d�:�Q�b`J(���8�K�����YB�w]�`����N��,qN�t�g�:���r�`!M[]�5~~�30�;B����j0�����"ڏ�HG���0��5O��{��@U宍�űn�x��mD0PQ��3�P8�4c�-:�h���vb8�[ ϞbP3H�I.�#�"�N�焊�>T���y��#Ei/������2��sh'��@f���ώ��$4�����"+�*t_"��*�"v�q��_�2�SLa,��0��i��3o}�+�!�N`��+�Q�|�}�1��~-���C�2�����x*jg���$1��L�D����ԏ���r����0Y�G	:�4zi��I�\i�4L�6��̄l��v�' T�����Z��z�>ll}3����Xg�ބ8g�Ԫ��Ԁ�˽ 33"%�Μ-´�J����Kw�@�Jfŝk![�Yi-��=��x��j�$.$lz�	��73��>�w��{X:�l��F^'\%T!ro�d��:N��.�芜��d������;���r��at��^5#k*����/�c,���xKi.�U�$�`���2�a0���(�?�v�L�:���pm	18Bf?b c���6hU�{�xrh>$�e��h�N�Yx���Ua���j���@-(pc䲖 W	x��_�([�x��ɯ�k�����b-)��@eI�����Y�Ѳ��g{,v����ڴ�L���׈l/����؃5����#j���|��#�7+:��_`o?��GR��R�9�{4t�aö��B��@�ܭ�Z=��7R	\A�h��
�=�N$�JaO+:���ɵ���z������hM�J���?�*����Qy`auE"�%�r�t����"��"��#������DX�\[�A���ZK��d�k��!�m��C��V[�YzzlE��0;Z���]}_��4��w?`���r�N���%�,�G�:졶YQ�_�
hރ=��%ASԷq@��Q������\���貘w��q'��2+g���]|Z�U���^���I�����B}�Gy`x��Եn��#��Tv��On���n��`�˵-���M[�M�!Ҝ��X>�sL���`a�W�;����pm�д��ۙ�椿��ǝ�.��:�q�c1����b���C�Z��Y�Z������:�|W���_��wq>(�W�S�<H�'�K���	���Ǭ'�oo$��P$6�Sv{o���jY�r��#���1|�2;Ȋ�4g6b`����t(d�,6iٍ('�z=!�B�Żh�46�ܢ���f71*��$N����+�U��~J�l�S�7c�4���:�,,�xVk���	�Z�?0��B7��C~6f��N0C��1F�W�hw��pJ6�{A�߀��+��5}�B��W��Zw?�E�;V9���;�H+�� G�K�@����v��e�̕�ݢu�M��6�P��	���Ng�xN��u�H����`���E�IS��\U����Nc�T���H���^�q�Iv�8�N8$�|�����L3���֡ 0�$��F��7U����5�8�)�'pװ�a� Nd2�5+�[\f>��n�B���jV�M�������z�[|���.��g��.5 �j���b��N�P�~���(�u���"t}�v����ku��������V1I �_�}	Y��X:�Wn_���^��q=NT�.I�[e��Q����,	OXp*@RW�	ȕ����f���s��疹�L�5	
��x�	*q�C��v���4ᶎ�)��H;�s�rRX^����э�p���	C����5�]m�h�1&�,;	o-O�EQaܳ�.�G��NX(f{��~5Fdj]�!=�h���k.E���^9H�6V��e��g!�k�\T�ΆИ/�'u�R\�Uf�l����B���x$��3t���5�D0��ʖ�Qq�7���z���N1|�q[,d	F����L��0/$�e�̈�=N̂wH[� �qV��dj'����B�ᖕg�}����������6�z� lJ���3���1�LŎA��a�J���(|r�N�:�LM��[Ӥ���-�|�j2<X��<��BQ2c���<��ށ۬�p��^47��XJC�ɳhS��Z5�pjY#�]��?�F�eB�|rŨ-=-L�x�SMDX$��_r~����_��oa�Gܶ���9Y�Ї-�@=�9e�)N�9B��0���%�0rK���`Dǻ����@+<�����r�F�)e};sA�Sh�G��� �;ϯ��̤�*k/�M��:\&G$@;x�J^�=�V���i`h�5¾d�/'mk�)�܇sv��ԛo@~`@0��ܱ�䌬�c�q?ܡ���T���A+���F�\�.�@�PX'���K��&��}��e���<&��I���N@3Zݜ��'oB����e/�o�s�N�q����+i��LF�k��qP ml2�|�Cr�߯�D�;�G��}�g11��I���i��l����s�� ��wr�Rl�q�K5�����ێ�^�3 ?ot�V ����`D�*^�M�q�҈��P����t��_,��\.䁴���ð�`χ+gG�Z�w�(���Y(��Y.�^�G抱�P�uv��B ��� ��W�k��T$D2f#���`�<�J��f��-����!��g�h⦡^���~�/	���@�3s����z�����4��\�ru9r����c�H��גna"r�y��6>ٽG���w ��Ö��sL@�����������JE_t� K��\��~�������_�+���F�+@���y�;j6��\%�A�rP�	s�P�٩P[������_ֻ{$��=��4�[nFE���>�����;�	����V���M,ߜ��Y��"�^vW�����&�� �3y|��9�1"#C��yƌ�Lm�^O���~�y���4�ݯ�2$��\��E�aگ�5f�eۺ�R$)$��_�g���v0E��v@n+�ʑiax��M��4���O�}8
�K��	��7���a���JtR$�_��~]���L��h��G�\c�w.���Q��}��ܥ�iI���A�ә)mG�3v�)�~�P���f��ؓX�}Zs<��ZY�1Z��
��~咬ww~�c���?T@c7��=��j���ɮj�sn�y!g�7,��2I�ፌ�RO e�W��'���Mǐ�	����XC(j�KL �j�I��3�����L��4��O��'�r/�ЅE؀�`�'����NZ���Y%�Ğ]c%�rH�p�~�?;���>��+�O�;�w�gT{��1.��������оS��� �d.��9�����8�M�FE�$	�Fz�
8A�Y�]�eֈ��B3�{���z�:4M6r���D���tM���&�����{y*A�Zڬ2���(=x��oy��<�>�T��0zH\�	��[���Y'kAR��R�:u����+�ɞ�B�R,,q��2.����=#�{]
d��,rD������6�"��I|č1kC2Z����!
T�&�X��/�f��<fܪ� T�F���1dN�����I��t��ׅ�|�3��i��&�D1��͡߇��M������J���*�!�2pꪝ�%|���}e��v���B����ص/4>9g����ƶh#���S��f�j՜�|g6#���)_���O��dU{a2m������!�$L��M(�|�/.�O R!Zbo{`j�W٥��h/��ț�\�X�9�M<�pk�'?X���:���QO\���2��۷���7F ��� ���H�28T{�9&�H�>8�K�QX�[?&��Qb%ɓ�1M���N"f�;sw���_����U_i���o�E��&�6�SVK,�EJq�q��}d�/�|l�Y>$F����gV�JDsy/�+$��W��ق���*vqB����y��%�MS�p��0��9��v#�k?d��K+J� Kiau�?�k���A�u��}x�X��{]'�g%0��h����C#��(�T"�p�^w�n�ugA��.��ҙ���Xg[�M��h�r�b�[�v��%�ĵ�*JC@����h�zq�E�w)��]Ǝ�H��p�mf��xq=�A:H����JoV�*���kT��Al��-�B���_,�,V#�>�X0��`����y-q���=��q��Jмش`�v^�s8#{��\�6�5�vVa1��j�FG~���'n���x>���q��3h.ԗ�Qݼ��.��[�Gjo^ ℰ���D#I�A�������F�Q�FC0�qScr��3�^L8��:��qԣčyv����H=��n�VXD�О�Xp�\���">4��ɘe_�,���1?
J�ۥmm�{X֪J�$C$ ��+b&h�T�On�(c��Sy�LC������γY��R#d0��L]@p��S$�z]��v6�Ԧ��+뭼��g�~�bob�q���"G6r�I����N�%��=y Z���w�r�0�	G�r�H�����l劸����h>� P=��\cdu�xl�(�Ӎ^x�8ґ��J�3��ReQ�#����̕�^w:͏��RXh�����2�Ar.���N�ǒ��ḣ��q^ ���|͖U��+:�+tNɆ�"-�6�$��~!{"���P���&$��ٙ"���@(��y��V�\B�0T��D�,�Al�Τ;�f��2����޶��͖t�_`Dj5tp"%�YO�i?D��M�aZ%@Syȶ\��m|UNhN:�� n�+¶lL1��a�ʐ���'�_��lcmaF?�� vCgt��kM�H+�J)ٖ��U�/��ô�DV���Xg�ڏ���`d�k4��6����	�ĀKIh�J�eF�p{,T�A���]Aa����?�*���u�}�*Cp�%��$��Ӎ{�F=HH�!n�8o�� {�nM��B6v弋�Y����? \}!���m	dѻ�$b9��:��׸��-�Y��B�����+4�lFҳ���j�t�CA��~�U즪���ag��	���Su[�OUIZ�p �W�κ���>�b��A�<�DͶ����"�%u}ONkL��o-B�ո���1I��J`�I���r�=j����'�����>p{�Q�<9���{�~n�$(w@1�����SѮ녎�h�]rCO��lPh!��j�������v.�f�;�:y�$�O9L�E](U�9EZ\�tQ���x�����
�!���g�w˼��И*q�GG���G�Pu�!�p����]�"�Q�g\=o|�e<Q+�&��?џ3���q}��qyS��{��d����H�(]�P�uK_#�����Xә(��b�g�����U�_*�I1�%���c(�B)�$Y�IZQ����B�Dc�h켴Hڤ����^���~�0��Q��5����}�x�3ϕȳ�q�m�7,�IA���/��k��+L�V�<�i	0
VA~"���v�1���h�Dq_�W�삽�~�>�%z�e0�Y!�Z�P٫����)�_B�zI�Zv+���vJ�C�U�����͵���l�a��U�ܔ��$(7�Uı�=y�IR3�X|�9�G�F�aȓ(��Z�79��K�<�T�<��n��9�����1�k����v��9#dp�^lD.�n"�Mtj�d{�a^�d�\JnQT���>�=�[_<l>�x��ӓG3��Xo>@����B>F�`�P�/;�6�{�l�EB �2wYϪ|�YZQI�a8KC�+����x���Ї֘ex��p��ೱ��.��E
jX�.�[xcs[�&N^��(�ŀ���F܎��	�w�𙽭@3�^�6��F��Y>���OE���9$�b�_�q���z�0,����F�С�,�`�g�7�����SdX�W��#�Uc4iˑ�௸��Ţ�-���G����^�rK �^$���~���;w3];��y�v���nDp``��m�I�P���&+&J��Vڎ��n]ʬ��"���aɵa
Z�\�����^�M��H���&�W��^��0֎�Q�>�c8'lgZL����4�حn�6���j�6�,��Kࡔ-8;���7�.��!��}�._`�7x��c�����GU}@��h8N��f�U��5��Bѵ����	~>��6|��Te�O��|�0�m`�*��D��u��^��!��\���'B��|Ջ��ya�h9A�_8�R����͊e\n}�`Ų@|���q��u/�x�����{vE2' oz�Dt�?Q��rۥ��Sbn]�«�$Bë�2E�}7����ѵv�I.cׅ�,�$��5�k�qV�{EkL�������u���.ʔ��3�>� �X'�m�~����K�a��oY�8���L�{p�����(|��:'/n�#��V�4X���Lz�P�v��%���\���T��^.��}&+���Pyq#��DP$��� ��8*ɳS�a�z�E�$�K�'��iq�L:�yE��YL�`C�J˶ś��LziiJ��g�]e%f1�3?f���sg�=	��+�չ���%*�A%���G�K�X���n����i��!�h�`�<��^0�W>:`Ɖ�E�t4R�5�!���"�.s�x�ȳ��lU�#�g�xx���ADI�u�ы[�}�)���cK������9J����Zx�X{\Y�(��E�g_$����E�2G�wuuH�Ѓ�^��2 ��̯����o�K<�6q���ҽ+\Ґ������3�)'�e��HQ�X9���Dp�
y�.r�gg�.���91BX��h��.��2�m�5�q�h�,��j�<A�P�u�\«�~�gW#�pj��?C=�P�D���^ �+�C��^��n�s����	(�8A=a�F[o��xZHZv����-<(�����p�Z�3vS�����HŽ�}�({�x����XN�pv1{��w7��������b��CrқF�x+h�b.�o�D��M���4 �z���u7�Jx>;�2X'���}����9�X����&��S2D�̡ b&ِ���<�J(�ܣ��l����j�C|R�@UI��gT_(m��T���UL$���"s#�_�M�3��ܚl4�^(�qZ���񱻓@�x�y�,����bY���A}9�)��s��
�Zzc�ښ8����qM��K�%=p�,�Q|�F��3��4u�R��h`�)�g�#t��D�ר��fK��d�'F_��DG��j��B�,����B��
�$}p�^os=����wf�*��6z��4��;� �1XV��~ �N�$�=�6}����ϬjF�/��v��8��SOK)��GG�k�s:��J;"XWG�PC��B]`�ʝ���{��x���un��-��8mŎ1G�%��w*�A͐�.� .��I\�B�p���M�w��^^�\�q�����썘(��F��f�3���Ս5X��s��]9��M��'2�(\�vWA���I��C|,%�l%\�᠄��R#R^I�ug5�T#���I~�4�Sb�����O���b�*���ҵMS��pX�g�d��z�O������8�͹�zT�d=�Gl\R^mS0�Vn@���<{p\�:��c�����d���H�<���ɳ]^���IKY���2c'��a�S꤁��� ��i&\��M�~���:>�l�[{F�^<�χX4��$�U,}:0T����X�$�E��=�K�WmI��04b���?�*5��i� 職�����=���k��m��]5���GA�QV���DI�4 �!߁�+6O��\H'�Q�d,��`��hd��g�5��C�gva��Vkp����l�iGǭ>9H4jF��$���X�R���D( ���w2~_��9�G9FH�ؖץ�����~V/j����p迲����i�=���X?e��BȲ��,�
���m����um��dN��Ӥ��|+��.�բ]�l�v�����{=��N�"k1pF�8����&���@�ƋG*��T����Q��橢(�|t+ �9�c��z_�M����1��L���n����� ֽD���V�w�Z+\��n��^�$�$8$�H��N��Bq���>�rY�a]\u�]��w����)�H��؃uAP�b�Bآ���Q=�����φ�H컊�x/w��[�aN]���%3�"~��� C�l\@�*���C|�"�t��B�Nv�k #jw �J/�#�c�oO�߸��3�}������#�[�&�K��[��x0�M���"W�6��� f���uA�T��W�nq;_<sb�j����!'||)`hҿϠOv������m�U���6F �����?݆�q�גT�!�.�ٯ0-c��^Z�knqGn^A��Ѥ
Ø���D�� 9�/�\L�x÷�A�_	���J����z�8Kܡ������Y�7�:c�c2�-a L�)�
����cU��9�����Nz��|���xI:O�<㾄ג>�kq�#Sfy{�'@��Z<�e�AEͰ��sg��v0U�E68�,M[r'�u�dP�-�W����j;yi|c���|�PU�Ĺ���HT=}����p��A�1~����}U��d�c|�K�e�5��O�,�Ԣl�eD�^a��+¢Kq�^?C���o����Q�!�X�M��l�M�!�b�6�M�s�5�'�=s�T��?�ڴ�kb����5{왑�5�n߸Լ��+�58^�b9ؓ����@{��3/6����g��+1�V�X�Ic�FY�%q+Ә�W=R��km}�@��%�����`֨%�T 8�3�� 	9U4&�eS}}M�v[K��6��@�quB=��ȓ��>f��YƵ�O���z�مkp�����l�m����^���O��?��~K	cٟ7.e=ΐ{��lN2+�Iv���FdW���e�v(	XZzR���\ 4�B�ल����1-�i*�Ӏ�U�\�s]IB�B�Z挲{ �*����mSM�� k57�l>Z�g��z��S��K<�]j
pW�$N��#�B]a3���)f	#G*��>�rr*��*��;����Z9>�Fl��]*���2�u#�-�Qփ�Xz���n��q�t�2j�`�,��g�Sx`A�(�+B�(PZ��h�t�<�^)m�u1�h��59�X@"�e�T��z#5�D;��@ay��Yș/���А��#`Z�Eb��h����2$)�J��1�*d�>~}��+ |�p��F����������fgc��-���ˬ���g �i�g����0s��?ő[R��tx1�-nC���T{W��FsdD�r��)�������,�a�!�����$I���sa�-����ea�x�%|k���`�������V�ԉ��b��.���a~��Lp�R˜�#���1�0$��@�Pܤq�_v��|�`c�����1T�'�T�bw�Q���XJlP>���6"��@PAّM/���q��)FG��8�U>B�������H� ,���-���J}(�8JM9Ө���H�& ;U1\' r�
R�F�(-����(ŵI>c���I�N�~�:^UL��֨[J �?�Lm���0ؠ9�l�@�=Z�������˫�2^���f\��lh{A{9u�:Έ�,�h�ޅ��T\�3��s>b&��?R�4 �1�M���FX�R���*����K�Fqɟ#h��iŇd�T�c ���V��*d)\P���S
a �E�v^�G�L��O�Q�ȯ�b-�PT{�W {>���a�bW�/Hu���Ls4��K9�@V��? ��?-y�޺;�8\��*�^���~�l=C4J��A��Y�81S�"���@Hϭ�a(ēX���~}fW�6�ۙ�iw��y��K��6��:��Y6fY\rx�A�k�Rp��Dhĸ|O1�!L[�=���%Y/���(I�&��7D��������
��O�Ņ{�ۥ��9��a�#\#�@l�||�\5�њ�QyZ��﫟���f�o���/�� ��cL�5-������W��Y��o��B���t�?����\�$;d&E���ֲd�o{����M�"E�������x��_���{.���􇓫O�,�����05�E;���,
-L{Lm�\��׍�y	ێ\Y�4c�d������k䉭CF&9�hG}IF��lVs(��B��p�$%k?X�����u*����e12��e��S�?ŏ�����EO[�vs���4�(9�n��s�]�����5u����v�Bl��G(2�j�_�� ��gw&�
�[gx �V؀�{+���J\&�2[�V����3�ͬU]p���0 T$��rPt�:BH��.�ݼ��1��\>�,2}�%@�A���+����EfS!��P�������3��T!ڨ����8g�wvǨ�W��0�2O�ՊU��C.7���;G�f�AeIy�-M���������캦c?Ј֘�[�`��<����yy�*�0O��1 ��	��9ĽE/����8ݷ[��YF$���[�ٸg��EY���J.��4�\p���T�v\�S��ݕ.˖?u8 p�F��g�9�Q\T�+Y*��ü˻�N(���N�C�D�<��J
�7�NF�$�?���⺲�o��W��^
[��;����3е�kz���@��ls���E0�C �Y3r��G·Q�ң9�?���,/��p��rt��G4�]u������2`�G���Z��Wh1�� rJih�/a�����ܢ�``�0�v�wd\5wus�2Ӝ?��� �6J��IӮ��,;)&�G`���|O�o���zIՙ�����!{c)�!��ZL�0#�p���o\f=�rߡe��=��u�RO����]t�Z���rh��������ǈ4t�[`�N<��yC�Y)�_b@D��}���54��
�!�ܬfn�UK�]{��(� ��a^�lRp����Y%�J�5m�γ�!�������g<������X#�З������3��X�&��˪p,��me1�"�|�Q�1c*��V~�==�z'{�N�7,����sl��ݷ8�A$7��(��煊M�h ��?ɍdh��/
=1'ĺ�|��~<�Еu+b����]J��3/0iy,����c<���W��V�B�I����06���Q�΀��ۻ58N���΋Sz�n	�s�3,�-���@y�D��^vs-�V���dz����4�d�U4Oa�><�/#:S�1�S�A+&C���0*�#��r��K�
�\��#�p���Ux��tF��������ش��{Y��#�ߤ��&Gv�Z�M�Nr�Ĝ$#��9 �A�i2Ӱ*�t��4�&/�� ��/�UG��0;?�O����M�]�H@=��_{ܵT?a�6���+�?'��E��iq=�EǮO��/G:�*:�������z�	W���$�O@�$�E���o�h���`̢�R)�8�R��Q
�խ��tE�˿w�9^��o�PRR�4g/��X�]��g_ǜK��q4t��8P(�xȈ)\7�>�����C-e]NȈ�����w�w��ȡ، ub�Xb.S�����1����z�3�o�y�o ~������o��Y��ޤ`=��� (���j��vp&��;ZBG��
���J_p��Vr�a�"@��4>�����(g\ �UeZ�JeF�e��T�:��qpr�}��N,��w��TQ��ҩ.��(KI76YI2k���h=��gk���˪.f�ʁ3��Ygmk�`n����݂W�OtƦ �4��u!S�$� G.�"���	t���$4Nr��a�(u��S7AE6�_1�*��Žʒ�,~\��T�^9��gvpqb���J�` BZ��m��.`~C���m8�]MU���|����*r =���^n��o�(G�_I�5�*}�NҩZ����L?��s$�M�
��1���*P�M(��w�a��� �6�����50���G��bq�L^<9��@U�Ϻ�|5�ZBŌ�~�m|����:E�|y
��150_6��*w�`U>���$N�$N��3�gD1��.�؈�4y�Sm6��_���/�m!��c��Ҵ
�Wӫ�n;���wB�_��,��[����G�e��j2����u�k
��ʳK\��6��a��	����?�h�a�oD��f� F�H�59y��BoB��WO1����'��WI�t%�6��:�(�Dm&]@p�H/���}F;w.^K��Vo�R��/r��h�`��;1!��Ғ%�(ϊ����EB�g�D`��,$�Ɓ�����6)���V<�=�ei� �CQ�P���Dbdۦ�{5 ��.�h�����#�͈,�<2�׵��8�M�I�����S�pR۴Q��U�B��F)|�0���'�S���ﭳY��f�B�BM{V�lSU�RDcl.���S����7����3��Et\�M��5p�#��4[�/�����0!K�;��6�Y��k����9���d-+�Ν���hX�"�o_7U��+a=Y_A�	�Iʒ����e�FQ��ni��ٙ	��$�Q�5�(f�v�B;��#ut���-��(��(%�(Hw7T�{�(?=埣6a����y@����w���w�2^ށq�xWV>���Uӛ|G-D�#���\�n}�<J`V�ʉy���ǡS��C��ewa0�̿
��|��e�w
�P������}�)���?��������zu�0|�6���SB4�0Q��B��������7�Ǆ����jw���' ^�
e�X s�q��#<� �a2����� ��3'�H7P6�O H2�l�n�3�Q��@�&S#g����}+Y�����w��t�"��5��=�I��*��9 ���P����N�������S�d��ֵ�r��\19��TG<M�!�D��p^u�Bす�,S����L64�`��@q5&�ቭ�<�c�Njvwz�x���{�>a��cH�0�M���%��L7�`��g�qE��l�>�h>�2
�G���ʈ)ק~��u+NZbћ[�C�+��Qg���<A�ղ~Y�H+�?�fR���:FY�怈G�-In�Jb�ݡ^h[g�����K]&���A�>z02mH�Y��;j^�K�n��v�Yu���q�~؃6�eL�{.��c�f����4 S�8$2t�H��)�� ���
R���]�k\� ��?�<�cv�J{���t9yR$��8�����!f��N5@|J1����������}+��J fJ� bo���-[�NL�H۟��^��ɱo�����հ%�`x������Z�z����V�Ķ>��J� �%�3�M�TE�h�L�1:��Gv%3	��+�ʰ��@�0�w�h�*'?߾�+5&��v���8n�9A[pVrฆr�l�_�u��]�I�7�ؿ8��,`Q�]���y�$�L��B�����ɆC	!��������v�G��;��,a齀nG+�+�,*p	ܺ�D�
ͶF� ���U(�<���a�;i�7T���U	�����ز'U��=��R�'�<]�9W�����$��� �nסb�~����X��3���~�<�Qcy/�$HG^�ܶQ�-��j�Y��n��{�r,o���%l�$Z�*cqX"�Łk��ם٪N�����v��1`��$]Є}�CW�8G"|{��y6Z��2<�*.��N���$IFI�z< sm�v�51	�R���3�ӽa�,Y�}d>I�f�[}��MQ/��2�-�f^�;�Lo��_�}lip�(Tɗv��v^u1�J���<�^r[��кl����5ٹ�!�x�2O���Dߒ�^��짧���ԒBiU��-�S�l�X��ȁ��m�yf�3 ���	n�]�$6"wù��p0R$�cN&6���I�g~qP$���$[�$	��q4��xw��)�0�ϕ2������ߙB�.-��b�}��f���T�w�<K�H���>˱����o�����'��Vi�1R��1�<7�}�V���RS��;�bBٯ���A-M?Nx<��'�Ux���յFM�w���n�cX��;���!5ĶQ)��\/��nb�eo�b/��_���;>>K��R4Ĭ��+�������]e=A<.����[�64Pj��K�>�X��ٖ���`[�P����-��JQ�vQ6/����s_0M�zM����P"?��=����׊Q�����mɮȩ+dM���?Ǡ�˰����U���z��Nc�R˭�|h!q�[*����fek,�MPu�p�.gCQ�|O�V��X�*�m��Կ5'�:�����D!|��o 7Hw�Jd$�KYl�P[h[�E�������k/��.}��f��ڐ�PY�&�(���_5�O_��	,�(��)����zf���)g)��uF���;<�����I6��&�9+�@�S�!pr��W�?X��̊�K��\�PW����{���=0��)`��W��c3���.���7�l6���|ɓ P�+p���Xa�h�~(��i���u��3�u�$:�0�ްީ}TsD*S,����FR�{T����N@����V]F�Wu��h�HSR��3g׶�*�#���O�Έ�J��8�7����Z��x�9��-H�+U����T��	��9��t�i�K�&h��O��\i����˷�1�@���<���9�|�خKt�77==�%��R�4dxhq���UE�UF�uf֢��l����ѥTe['݈dv����ٕї�P�C!�݁6b)T\��7�T����	�n�愷�`;����2�H/��=k���ǡ�C�QE�d>bsޢ�>P�L۷D��W�X�k��`n�\KPVn[e��ʐ-O���S	�E!��v�0�r���m'�z�v�y=�8r��U1{ǡl��p3��Y�h��t����Ϋ���קpB-
x�m��q�<�=*D޹���D��2�L�s ='��ʿ`��a�]����/���Ɠ��J�p7�(}Vl�A�T��_�p2�|F��dX	�n���O�.�Jݢ�8�sf�=H��n.�b��@�'�W�e�y�vc���}��P�6HH�>��2��[U�#�#l1g�>��%�@x���Y��}[T��w��w*UE'bG��۰x��>Uq���r�ؑ�~�Tl�Wy���D��J�עD����_�
cH��=�<3jC��)޴���zI��$>F��y@�"h�l[X[�j�"Adұ��0����n�R���o�;�	Ph��\�N<vS��(�yƶ{���op�N��w�����. ���:h�9A!��1�|<�L<\Ki��-ݬ�E�\��֠�z��'j�q���:�
�t;�B�8�\%S�C��ߴ��l��FS��o�ӠZ����9G��3N,R�%��2{������{kW&Z�Ŋk.BD���w�a����&�53��ʋ1-�=e��j5�>�ڪbN]���+R����N������9�����"��,�47� qt�|C66L~�+��0�N*"��l�+	�}@N��"IT˴�W��<��ft^ㄙ��NnTuI�N@w>DL7���
��F^r���D��;2B����C�������ϵK_.�fD�b���@�&C:a�"��(�Y�a��W��|B㪪�_
7�G����)�n�X��T#kO��i������O��$��f��^]��#�2T�q^���񄪁(����]�x�.�8����m�TM�����z�)M�����6��U����q����v���^��o�h�M� ~��qU���=�hb�<ZNF�w���`��9hĨ��D�sV��Vox��5& ٟvB"=3|:�ή!
��&���k=o�D6@����X��J��J�eO�Ɉ�aJ�uV�h�
�T���ܣ�j�O������یV��.�>s�(�<T�(B�?)g�P���������-��_n�b�G�hOo`���靟�����s��E�Жw�t�F�OJ@HƑ�@'��lHpdQ)ih�Dl����D�L�*t��i6 ��l"�V��9�ϵ��
oc��4,T.�l��"R^SVj���6*��UVi��ǕM0�������]�_ U	#���~�I��l�Ji-�ƈ�+e�v1���˚��UF.��!�S�mL1�벴��M�������s<�[�oQT"5{-���R)W����8�|�f�>r�v�z³C�g.G�3^�/�<7G�]��6!%cpԹ�l#����'?�Ũ�����{Q �>�y�ޡ~�9DJVmy��Q�u�T�n��p�B��~J�����}��T��T��9�ϧ�����Mq9� �8��x��yy����|�y(+�uC��ņ���-_���H���HQ���%�5���^N��Qr�mK4��S�{IY���h	I$�1���bEa,T�ҼR!Sfi�՟�*�,37�9����B���2��Z�n�in�$��=9��v��=�|Q�{Ī�K(�$���y}��c'�5G���cz�� �N�O�8vWO��<P���� ����2��y>�.�@������p��u�q�#��V�휗v�Y)��i�[P>�YF�@ 4��AD�*d�XggRi��A���r�p[
��4���o��"@һ��v��o�)�N�(ޠk3�:�P���$�]Uw/D�����J\�v�k��qV�i|��9%��u�� �Ϻڈ�C���}�̗�yV,����+����l��Z3�=�p,TGjxnw1�_k][k��βoaՙ��8l�c�n��4R%���ed�L6�sP1������}�!���`�:����]ܒ-q ��s�@�V2����[&j%���+n~�9]>a4n������)
�_ݎ[ �����]�vGgfu���� ^@J25rwJ�[��	����c�L���/�ۇ��A����?�A�a&�̰6xi��<K�V�@�%�H�u�&]Eq�4<�hJ�E31^lWC^�ۣh����7+�Wϝ�|f���_���4#d�We۶�o��n�k��`�gyO�Ef��vcm���\ѲlK΢���3J�B�>�&a�y���aE���W�~T��m����W�k!�l@	�n+���_�g���{��F�{k�zƮ�f����F�K�4�)"]�[L�����a2�p�6�އY<p��⁳�M\��I�"&</_I����i+Y@�P�q������<�zˈ� �@�K��c���A8��u�NS��ܞ�5`��]�#o��p�VP[�;�/�>J���N]�u����H��,~�ԕEj1�-a�%��R�-��=�yt�Xm����o��%���-��J��<'�#�x���qYݦ��W�F���4�#w�GZERNǘ�J$��/Xf�%J1� ;�b>���%��M��N1�c�9�qh�`?��O�.��:J�e1�(�E_�914G�v���r8�">��sQE��=K!����/�WI��U�Z|�F˵�	�f�`H�����	��ρ�g3��d�F�.J"��{���0QR-xWn��]n�\�'D85=�(]�q����w�
:��F\�Y�(=vQv��)K��Hb�]Z�E�K���7���B���",�����P��,�O|%s��.D�e'������۩��͈~ Z's�Cuc��uIC� �����9~Cx�s	ik�D�A	}�1]V���cQo����Eƥӳ�(���y9ʰ�!��w���`�tE�
Ѽ%�g��f83�6A##�|�,Ǎ#ɝ��7+�ܭ5��5�TF���O����@ n0yL��]������{����s3��6�5�;z�\�*U��q�����)I��RT?ԋ��}�=֪��6k�mb�Zf���<��Gv�5�����m��($���P�b�{(���HiXs�n)6գ��]9��bR� /�N��ю���_)��Y��
�c{��n4'���aP$�&I��FxT�)����5i]�r)qM�.}��g��*������Έ��(#:7��� J�`��@�^Nb���J����~:��BFj��:������J��	�4 �����i�0.a{���z������>�A���J�F0�L�2��n3%Fyi2/�U�y���=R�����}���O�@�5&�K�\�O�W�(VM@P`
s��I\�к ��*�����>�j�ż��������+1�-��El�uߏ1a���Y"�fl S�b�$�8N�;�z� ����r����-<�Ċm�S��]|?/G��Apܨ`o!D@�. ��}���(��kkԌ$ʧ�>otG&�E'RXnm�U6b�w��$����>� �J_q��AQ�<�+�r�DM$�r�F��mTp�ņ�Y��ʑbi9�T��u�)��xk
�:}�5 �<V%�w�m�+�t�d�>��s#Ѕc�N��s��y�3��)r���L� Ȃ�#���w�f�r��Z�aL	�����Q9��=���b�h���YL�O0ǃ���NN�'u*4>~g��4�OS�k.���h�3z�'s�M������#�%��L� ;���Àsg��C��v�68]�@�����F����rf�{�xa��;J��n��<�� �D����w?\�q��j�Y��l<!�u���,���\%��a#M8b�"�^j���G!2 aq |#헦��@<�*/�ր��:�n�&0��4ԬT�n�t֒{����k \'��m��R���	>���$B!�$i*n�C8�;9���l������V�A[v�&Wz�S8ʾu���1Wݶ |>|�Aq��5-��d����Vv��#e��$i�Ӈ����5[�l����#�k����!�諏_�}-�gV�hB���;�Z=_�- �&	l��̊5 ��ݮ�#iE��'�`rc���T�`wOyN��րC6|�\��xW]d��r�H��@�{��	��*����^w�
�r�%��S���uS<*��x�SLml  E["Ժ����>S���:�*��.�����X���:	&�������i��ObM)���)~�?`�Ns��A����cfq��|δ/�%{��&Ʉ��e<���bq4Mʄ��f�c��gH��b��H�Hԑ�Ř6U��#Y�V��@������������@�e��ac�-�7�jY^���^>�<�:�cP!��yv�-E�Y]<��ɼʨ̔��V����
�|���_G�g�%���fs'�~�~���?&���Ҹ����^v~���ŋG�)J4r�"�5��X1�h���å�@�����OLR�ն`��zp��"�ﯟ�b�+�P~�/��[8x����wf�8��"@�P2���S��� ���a�C$Қ�ľ�ɭ�E&�?���$�����r	w�F�w���FÔ��0e42��)˯>�m�u3�������>,��v�2zJ�)-��&����)1{o+f�a����ꪃ#AN������(�jgX�8�<0Ϫ=�]Ry��tY�*�N��mF�g.6�XV͛B�C-Y��l4�f���4��	����*��\�a/�WP��~Q.��I�;��@�~�(n�y4����iz��\+UJ�g���F��[q.��tr�AO�kQ��4�C��_�
�y���v�|���Ő�iJ��2���
��z�h�"�j�M��WsV9������"ſ���v���N!��C��D����z�8�~k���S�H��aO�MB�s*�
��ˏu�p�4_
q`�P�����A�J2���b,�>GLۑ\r絏bD`�+z��V�C<���`nc�M�����e΂E��,��!'섒���tr����m��f�?��~�!�⧑��Q�֛�W�y֞�8?������x2��E�0Eg&0�b��}��e6�P;�Rd�x6M]f��s��}�B.��U���U� jd��s�[۠��:��3�ˊ�s�p��w ���;ވ��ȟ���Okϟ{*+�U�zcQ��pk(BH5����'�:����?CZ�O�SW�m���G��h�E���g����c�.9�f2�ٙ���=�
+AY�J.��[���.� �q�w�7X��r[մ*�����(h�(���ŏ��`�rAk�.��=�;q%�C	�n΅����]�����~�ǹ���V�^3g���ݽF���J�87�8cDF�Lf*�=�l]��7ŏ�
s�ʥ�'78qВ���Z&F9�ȝ>��g���i��d�����'��B�nL��d��,���>�qS��c���-�
�ՙ;���`a�X��ehpk���/n��;<��?��H߈G���,PTX �Ҋ��/*w�H�|����`��$\q��mHPx���H �"��T��6�-��B}Ud�;��w�Ƀ�ԝY$b�t�����I�T;fx��e��ؐb�� àp����0M�U�HN����I������W8�6��O��f6޵n^B���L*�bK8��$���*AS�ѣ{ڸ탎nN��[��r:̼�� Qp_f���[ŕ����G�!i�z7(F�>�ŷ��}��<qSdԐ�FF��u��mI��X�D��m��J�J|���4���5n��H�ѡ�7%��L)�ۆ�z4��^9Ჭ7�J��xs��?Yg��Π�(F�y%/�Aj��ڇW��̱9*�K�pʙ�q�L��[���{��4U�t=$�(z��h���j�K����ܳ�u[�A����%o��܈��W�LȀ��	~�ލФ�x'��h��d���ݩC� �<����{g�*Kt_���t��K�UW.��J�]ʾ��"��@tѐx�xR����8U_�����#�@ @�k[_Y0��[����z�ʍӵ$)���f��W��B�W�b���&�R&;��覊r�@��d���O��+D�R�S��ơFƜyR�k���E��g�S��
�#��9T�a%�N5\������y�U����sq�P��C	ֲ�t,s*���������)���P�KQ�,��C��$߮Q�܌��5���츊n㤌�=�:U��
y��H�	��
�L ~������[����2���h�H�$��!�� _��.?�\�O�%y3���������=M2�:�v%%��xP@`3�(��>�2g���,1>�h�ߛZ=T�?�5��zbO�}-'1������Σ��ӭ��tޣ� �X�z�^+=��Q�H z>���)�j����+^�\�6wd:��C�=d4,�1UԟL�TK��1�%�jC��R㟾�#�~bV%�c�̾��av��鷞sP^�3�{B��]�r5�(}�S;-�d�/qJ�l^`+Z��~˰����J�
��k\�
,Kz��A���": �e� �4.��mG.u�?�w�؊'�h�E�҉	�*++#��E
�l��_ꎝV�����|� �o�Q����c0zRC�E#�4��T��o�С�"rW��#�i�t��T5t����`\A��?����0��ws@\�q����|G#"�Z���`��I6�_�A޵=s���/Ө�,�����c��1�`�>�|��(7�k�&G��R�z�sz����s��
��ĥ���8a�*�����\2���Ϻm�/I�d���f�y��?0�qq�29Ie�)[ ��q�����)���Dnϔ��ʇ �x�ixL5����p����6��`�Ϟ����G�P��UrC|��;�V1�w`�h��Hgr����̺�#o��3�Ϳ����@G���Ԃ��i�CK$���I'ī��;*0P_l
� dݒ�ʼ�_tF��oꌴ���U����<��}~�����~�^+\�Qy��u?�+wjw���p�,��|v���R�D^ze.�?Xux����(!	����Dc����Ɲ��1y7��l4�!��{9�6Z,�e�?
�M� �|[���,Ҁ�u�J#�ۀ��-�@�u��"H�7�1?�x�,c9=����u�/�������B�'!
&����K4P�LF+̝ �K��r����4�{)�J[�(T�"�wu��Ⱦ���fh �;4":���`�j:�*-8+�ˎ���v�ɣ�������yҏ�R�8���*b���*�P���~���8��t��� L�D��_��'eA�<%�`�Q�gʥI�qc��Q>�~�f��S`!h5�FfA��6����1m ����p;©�`+�bN*zon1U�O������{+����V
���6:�.��۾�X���5s�t
���G�H=|���v;�k�p12��k8MJ�ɤ�<J��Հמ��u�xl�p��&��t�v2H�0F4�ƸlưL4��m��BU����s����@'0=h� :�z���\��p�|�n6N)�4��E�%�H��_jeþf�����:0��_�@h^eE��R��Gg���0rtBsE&w=j��m�oR�ٟ����FXP&31�4�'ݖ��SVl�i����d�uf�G�(b֩�{y8��FR�\�p� 7[�'7�摒���~�Rk�0n�4�,���&h��d�g?92
3��8A��r��U "^g�/�>�MA[�v�@]�|;a5M=GJ������d�[�a�}�e��A�
a^?������p����)T��ip�������̓�1�w�'@�����%}�I�{�8l딺�'dz���4	���:`��ۗ׻uD"��b��'`y��CG$@�>����U��.�j��h�+؛=�	��1L�q�5)�P�4�,�](��`9�C�z4�����i0���������pm�[V��殌�C:�9�H�i�ӖlL��k�� ��Q��uk��B_)���R� �͈�	�� qdҍ��ؒ�Ƨ�N��g#��%���m��<�:��L#TM�QjU���3����4ce�m��:�����K{�*����,{�����V��܁P��'�X&�1z `㱴W
GK�6�M ��+�� ��#�ni��Y��������4��<ͺ�+n��XBL�~��F�f@K��]���*,}b�^-&����9��AV��7�L@2BX�ك_��e`D�����	`�i��@α^�dEvǏi��l��aS:@��_�>�D�d�P0��j��ywj,Tk@�f�"x��1b��Ʉߌ���_r�͔6����]j� ��e�M����jP�, P�Y��+�i�~�v�:(m���5�o�}ѺY��)1(��f��zQ�>t)bd<���͞�Go�N��"����k)� ��UV.�v��
H�6�z�(��kj�nMЗW�h�'�>���g��$��n8�����*4�g��歧�xS�6� �ኦ�vGǑ�]'�;�?[!�x�.�g����xj
�������u0��j`m/�e5��BS`�o��-g�(O��M�w(�3s4+V^��Aϵ�ϊ���#��bX�A��S�SƏ���Ө����d��"=���SZg�0�d��){3^v��f~(Z�M�iOm�)��~1<>�.����Ys�59��d��}��y��UCl�,�)��;C�&T����<("���+�f�x�R;S�t�EЂ���SQ�=�r�rܚ�*Lg��bzWj;�4*UV��I�J�p̐���v(���i1����l-�z���T	9B���һf�$�L7�'�S��r�^����r��$�|�sZ������KL�̜E%�����s���w)rWqH�5^a��@ڷ������rU��*����8�`�vřs��M�,:>es����g�	�	��u��Ჹ�^ܠŨ���K{�)���`���>������e]�1�����j�{NWH��]0�ѧ��[�\��W5\'�Q�9��8i�[s�?p�%~\yD�Q�	������%U�޶��4#�d�s���@uw��ּwCk3׎C����'Ш6)w"�\�n��iȬr�]�}BlVmɽ�~.�
�J������V�<�d�K��D��m���R��0��M3@ӱT��}��C��#K+�30��O�z�x	ҽ���9�&�6 �l۴��>I��dpޭ�;�Backf*�a,&��D��"X�F��H%4���,��%(��OS�(��G�ș7�ﲐ�=��]�����3��V2o���V�|�`�Y��W�,�dKĔ��t�8��ODGK˰ԙ��@�2���/��AW��U��Ȭ�5���?��;|�r��,d�d�9�����I�SB�~��F�{�Iܶ�P��]���t����7i�ȵ>'9���e�Z�?u(�V��g� ��j�j�Ji��c����Ķ�	�]��Q�i'�j�hZ3҅�۱<$A�X���Mܳ��]Ń$_����8� ��?c~ް^8�P,��;�gevG2�Q����+I�ß���گ���I�Tm'��mz�k�ǌT��O��8ʮ���nY�p�+E�U�zn2;��T�~��	�1������M�OԮ�f%ge�(SL�^^p�5�qO�xkѬ�p��6d�\zք����6�zj���2�1
 ϗ��l5��8�B>"�_ч�M%�Lm������!�v������/�Jz$@a����}^gC����>ؗ�bF�y�L;���khyV#�1VP_`s��X��"Gήz�dk:�|z�8�=
r�����wimU6�g�P���X�Y"�d�6|OUD�$��q,�S� siV|r'�����W���I��o!jj�&M���Rީ�/DӟA]$콰U�%��%V�z�[�8�p'Z>C2�!�����o)7m��R��q�ҵE��viY|�I�u�*�zCD�k8�%�SZ���v��|�LW���◩�Y�R(]7#��vݜ�3 V��墥
��4o�%�"��\��HP� �]�mR)̀<�gաs+����0�J �U�q=,-�C<��Ǎ:�c�(�ϾM�t��)0�yŚ�ax}ܫ��4�R����~_��z\8���	ƕ��hY]��C��0�ݑI� �e�LP�UKS'�m��d���������JE�vq�*\����٤�zj7ó�`��I%���p\���JeV��֧B�Ta�['�c3����;�q�vy$���C��_�`�f���2�|18��0�[h�QF���%#e����MDr�!��j�y_h�@��@H��N��IH�;]bbh��H�@�I�)��hQ��2��Bb�﨟j�ݩv��<����j2�sA�������Ƹ�'����/�dq�����u����F���浃uOe.f���_ �;�h��^yױy���Z4'�z%l#3ЉB0���Le��d.�>\��b:pA0N�ë���j�����B�BЊ5��h=1>�3@t{��fm���J{���B�O���pkN�}��H�8z�[��n^�,�m3k�`��Ǫ�
����3�]&7��8�1�"<F�0�㢸��AcZ_�?����L0��{|�w���V�)H,-Z��K巫H?"���ޤG��n�k3bȖR�eP�#S���o��}��+��8|s�7������bR�$q�c�3zDW4#��I�>=+Fq02h�P[� �AsyB�d���e���Cn(.Bŷ�5�r8����F����c2�
2nߒ�=��@M]��QR[至Iy��Li��`�@��陎hͫ�8���*)	���m������:��ņr��M�0���7Ribd��� ~�e������Qz���3�no,�j'p�w �Ե�}3k7W��+mG�CϘ�����#⭭�+���D6�=U��Y��d
�.7i�RT����OyW��Z�Z��4)+KΙB��"GS�$@q�L,/�R�>�s�t
p�тr�FN���o�Q[�f2֒35�k�5�~����Z[4��>�уd��4��#��0���4���t���2'B��#[�˟v�s�+a��P�/���Jfd��8�P.�>n�lh�͗�*��HA�-;����~ˋ��O+8@p����Z*�T�%Z��������,Kx����̂4��` ;h�F���x������ �ӞJ�fR��f���;T�a���˪���G�eO)@DZH�9����9>�����k��i��ڎFrq��Q�B�3�����Hc'��Z� ��*��
�����InL�E�O!_�9Z�U�L����TW�����Ф�0>^���!�Q	7�7E0c������ 2g��;Eo�Py�s����bջ�$^?|`QT�wfs!�atK7�\#��~���Ic@��U�N�~4���0B��<�w>�E��3w@?_�
�fA��\M��<�#�|���&�f�$�Dc+�Ws+�}�8����P����8���V��kg��2��
�+�W�wɿ}W��d�zp|�->��7���)zGEamU�=��e%8w&
ccPV�����{�i�j7�L�T�림�ϼ�Q���!�I��@��+�����5Gw��R��͋��M�ݡr�	g�i�;9��"�<DP,ykKV�2��1_�g��)���ff*5c�S�Ʈǌ�@fk�[�D5s�w���#�*�!�"庂(Pwy2�dt��#���=Y���P�Ͳ�P �a��l���#9�e���@�8�`n 2����T1���!��+�
�pi�Y��Rֈq�`���s]7�&�b�QD��E2U��_��՞���+��9��]?,$u-��ɗ��a���(�_s��\������d�H��χx\bmo�_�>�x
h������Z��s�e1"d�7UHL��j����z1�d���6%`�m
�@L\%W�R�{Si�Z�Fe�&͖��-|S��?-�|�Ȣ��y%��
��Q��v�X��'N<U��7�cY�����/=�q�ԪT��-�a�a��/�r��W���k�Q�r��݆Q	��9K6�@�h�����Mf{�ڮ�j���C�d����Q�q=��y� �.��9�c)��f���'Z,�u:&C)5�فy��>���6�������6�E��b��0�a�l�Q*�Y��3K3�=�'vQ��o@����E�^�DmR��J�e��1�#|�oр`?y����M2�6�w=+-χ�Y��,O%6hf���vȶܹ�R�=�M��~�/J?�#��*T���‴(m���m��j��Dw�쵤���/�z=G&k*���ߑ���Vѫ�2ͨ$�<9v:����O�2�fW]Efq,ܗ#��@�`@-/�K;�'�g�'�=/��������0�	�+�bn��ͮ�%�7��t��U�z��/#�8���?��w��Ж��yVC��-<,�m�q���h F[���_Ɏu?��/��J����tԚa�����ދ�%�Q���~av��JI2�r��;e�src�z��P�Jf��n�2�$$N�>���y���(g�a|س�zQt��l(kZUU�h
��FBlY��ٸ��*I1�Q �$�
	}A�a�\�	����? �o7 ���?�E�rv��X��r	f�n�VS��
�K���ںT�B`���k���I|GY�%��$vk�i(���?��I�-I^'(R[�\���I�芤=�
3����@�	�R�+�]���^�%�u�Ѯ�q�,����x�C�=	$S5�	��L�gJZ�53w����i�s,�ŉ����N�&2�N��j0����J�e4ZSw?�r��6�p�1FB��ʺ/J�(����]^a>��ʽ�����h�{��E�Sq�FQ�5�!BKrpCd8A{V� ��]���a�De�rs[�p�u���_��/�Ƃ�Z����.��&t�&���\y�^"C4��kc��`�F㊃�u��PQTu+�w��'� I!�����b�o& �Rؿo�X9�^�BpSu���YAˡ<���n�I�D�]m�7���;��m@��?�Fk���©5ǁ��gd�	�Cƿ�m�NNR�]���.�㝬-+��г�ص���ߢ�r�8G��Mu�z��xZ��	ǘ�z���G�w��S��I����R��Ǉ�����eK����Ab�Z��)�O�7G�U1���L*v#�8�� 9C�51��N���2������J�a�?�0�Kr5�L���?� ?o�?%	������F�"�R�d�$5�Q��īw�!٥����e �	��є�+���r3�l��t��h�,*0y�
��%����춄�F�+�H��9�y�����mԏ�k�j����޷�F��TM	�O�mQ��X�	)j{,)�ԜH�H��1�R4����J$��38����w��,<��+��	�UH��k�=�i�	>|'�	VS�'vn�XO1k7K���;�s�
�����l�6ii˶�g�	��<{�Ze���uFx�:�R^ǉH�_١��ʡ��A��I������u[��o�������cB�3 ��?)�b�7J����M�.Z�ڧ�O���T�m�M�"��o��?R��w�M��r`��J�o���t�����+j&������ ��a�.vZ}=�N�&��]�:ۑ&�a]�����6[Do;�cA"Y�}�:���=����J쐼����x�Z�nCս��8%�)��O;+E:a��3{8���!�,Sм��
� ("M0ŐC�2���B�F��j���n����
�� ��U�Y$\֢�x�hj�mi��%A�bm�}`�^o�*v��/��rAak�nW��XȦ�w�7y�!�=1��ݡ�o���=_��]�{@yn�>�4v|{��Yu���L1?�ý�j����n4{_^��2�0W>��ot%g�N
H�Ņ�����@���i�U������+͛�ڷ���ة͑B�3wwv4��\������� k?$�1���m�d�q�Ԗਸ਼6W/7����+��/��&H�=����B%���^n%'�3ҭH�.�O�E:9k�x��|�N�~e;�
���0)�]��}��I�����/EZ�#d�GoG8����!�vzʘ���r6�xSl��Ip�дV�L�Wflɘ�1�i/\��X�®0|4˞�rl��Ό0�
�Mԁo3~�,�4�@̵�ұ@����A��xP/gpK<��K����Go� "���%\��O��Q�9>HI)U �(��]t�-ݑM^}%�9	.��ԯu��<����.QBkc��+�ŵR��j��Ǆ7�rI�-t����V{ְ7�}��@�Wq��p����D��!
��%�P�R��:̽w�ƶ	,���uX�6�g�p�^Xf�2���e�[�ɾ�N9WB�Y��D�rCC7"/2�&�0��'�A��'��"�a��3a<��Ӟh~��$�b��{��U8�{}���`=�S^~��[�3�
PN�P1�$zN���J5��R��7^FYs���s�ե�dbd��k�I#D���=�T�N�z�,�͐G�7.|���ϯbQt"vj���Xhd�uc[��k^�?]�Ϝ�y�e�'wM�`�����>��O�ıH��eRoO��H��� ��j�x�蛏b^2����v+�T�����/��N���K�ތ]B�6�c����bf/�L��VC�i;ʣ?��=EP�|�u���t�m���"n���P�V$b�'��&Hh����m���a-Z�:y�9H�X��뜕�jgÂ�����I�x'���f������:f����ـg�a��U(�P��y��_��I�9��?Bs�J�HԈ�jߏ#8�a��X�4�M"��r{0���[��̔F��9h`�᱗��߆Z]�	���ޢ�����elM�TY�^/φ��h_ �v�(�d�딮�=��
�^���$Rф�!��<��R�8rj �rud���P��n�ޘt�M�n��T"�L#'�K�Y����((�o��5�)IQ��G'M�{����~]�<��v3M �U� ��됰���wd�]���0;;fK��M�V�\�	[b�J��$�0���N{��7`�A�B�B�_1:R�
�v[%g�u��D<����c�_��oq��<�9+���_�C9�b���r-��l��o�P���j<���������]N-��J�h��(�F�F�2hqKbI�yOP4{sW���(�j�,Z��V�w"vj�( �����;$Z]dޛ��_��ƴ�����~�����w\l�3������a�.�T��6(d���*��I�͚?R7��ڇY��b��
_�`��J;���ǏG�"��{�� �UYR��Q�	��3`O!�%�_���R0*�o@3A��ѱ��Dd�F�IiZ�ד�E��6��Xz� �K�[V��c�!Y&n?��@�G��E�Hl)1UAb�e4�K6Nvic�fw�6-�U�.�m�@����bDz�hsf<��H���tD�a�����fn����
����hm�(��A��!%F���t�cfE<�*��qC^@Qjv\����G�"c����P��dT3��%�bH؈&�r��'�tn��}>����*%4q��<�*BE�ת@?�����
4�"q����6B��5�'�JlU6�
ssG��?��${��I��/>)�2�t?(�� �U����G8xy�Ql���������"V4ǎ=r��)SOo�t�y��n����M��X�YoLoN�<fD%����K��e�/�qU!X��=ŨJDl���S6���&�#d��0���q5~+=��'	都~�P@�Qt��&���^>]+MU�5���$at�0�4\�������4�B� �yZ�n���#B�d���w/���i"o�J�%� �U~���\��������WdU����b�>��7�O�X�����Z3����Ӯ��3��}�8��!����K�S�6�*�=�%�AP�+�1ȶm����@xR�6adL�M���Gi�9�f�;Q�iIy�g�歜c�k�Ԃ??���� m�tM��l.�5R1������_8���������� &L��f%�`W��d_N��K/ ����{OȚN���:�6D�/ǰ��cj��T�H�o��R-��kb�f=&�%݌��q1�6��v.�lN��u~��0��?���a�%��|j��������l��f�H�]� M��'D��2��x6jD��i�����l{˝�w2�vK�43U �aupE	�}�TaD�^���� ��_g�o�O%������V�)�������s~�;���3��9�4���n�=����o�K�zZ8�.�,�u���!�|ş%J�����XN���c��6z{ZN�m�'-�O�w �O��uۥ��ٟ˸ƷLA�R��!�'���"!��u�:���YLz���"��\b���ΰ-�-�l5�y�0�Н)���c��{�h�)�.Sb�a�DJ�h����ClJO] hG�L�P�!�����{��g����6�nx+۳O�udO1cu���%��ƨg��w��ud�F�N�3�Q��˘��l��| �
<>}%!9��W�N�1ݱK���H��U��~}5�	�BH�0��t�N��t�a�}�RW<�OV�S�	Cf�ʗ���0��?���@�"
�����]�"�T�#a$� h�
�]�|j�a�m�֖s''�'ڴW������D-tm�͖���{���}���Lq���П��v]��5҉�C`U�>8��I'�w�i}w0���1L:���6�X#�	AmN����=d��C(� լ�V���������7'���' ?��a�u�J��#Q�	�Ǻ���e[/uhӊ�τ񠠂�q�!�b�$*��_�$1�Z����͚�&<O)=*y�^|��X1�������y����>�$��֝�[~�����[Y6eR��K�6M��]��[>�Uw�*�[�C�8�����Y!��X�����Dv�ių!��Q��>������#���.�y�%��ߕ��j���!�o�lS,�ww �l���$�}�4"�ῠ�ρ�#G���K+h��I����J��ė�2���-1p���~�F��W���\؍N�H�ݦ�^�Y7ԎQ|�m:�?Fw�שm:q1���:��{��S���~ӭ�`p�����m��; �\��M�"��7RU:�*e�p)�邓E�q��Wa�nh�]5�� 8݂S�� ��e��}-谻��F�i��ls�ū�C*wg7�'!e�C�ۼ��G�I��z��òW�׸}^��ݵ��lA+��KO(y��Ng���ӡ򍞟4��ڡx*'2��*��#���B��ǧڈ[y�����t*� ����G�߰g�Z��*5�-Z���8*�eBMp�S�{F��L���Ў�(S^�5.�"])��8p�-y�����&$h��� �$���&���®����8Ս(��*�X`�+~��tډS$����>�YN7
��R�JK;L��R�g>j��2�&�|�_L���@nH��(�`N2G�?��T��0XP�x�|���a��;{/�[.�q�!��ha�eP4��vIu��}�'�P0��@�؁���]���rw�<ζ�im4�W��g�Zs�z��U��4�dt120�b�y8��,H����L��Z��^v�����c^K�&������z�͸��q����׮]����t���n7NpV�2�j���(� ���/���'�.�����pM)S��S��;�!�D��pF�SY�!br��޲j��=��ڬ��3nҜ�ǜ�Z
ů���+x���rm2LҊ�'�N�|O�G.�oݑ��:�o���ؖp;��?�|{��N
�|�Η)�wz�ܔP�0M�s���}Xu�'�4^�tʬ�|����}�� ���;� `��+ãS7�9�:�Օ*�mk�p_�Pĭ���&�m�7���Xq��Wgۢnٗ�����pF���[y� I�Xڷ�l�E8(B#�%X�񽱴7�o�zj2G�뵉,��'��_���f�Ju�,�ã$,`T eFT뷀Z2�s�[�\�@�`2��n�,w2���
1�X��ph4L2��s��D 9��@��b�qu������$L}C��?+(ڈ��~%�,��,��Y�1DdF�p��]j��c:)S��J�������V�KkG��iF�	;	~S��u�$ ZR�vhѫ�K�3P�NC�������Q����EY����;�WfĤ\-�Py����s��
�Q��z茤b���)������*&KB�b�,�!��/���]��慐^�?��lo~-@{0���r>�:0	u!
Gnk'��;�%��R?C�|��S��K�2.�YQ6v>)�}���O9�J�f������n牕�7��2K+�ؼ�w1�Z��ʆ�u-S��ޫ�Ew��](�����z��0�Yf�����da>�أ��˛)Ly;�(�Fi�Rg�VX�/2��DK���nS�zR_Np����3�kh��Z�7'h}�e�r��R"o��8A$�t��Qav�_���_2��;�oG�&Qn'y�*�nض��b�.y�%�٫��OB6se��،��8Gr,��J+�N�r��h��k��|,O�%'<
��%�D4;�X�.�IEB��<Y�F���;?����nd?	u_I�k��?M�pvd=k&������~�Q,�ȥ4���������Uj�A�c�����Vvm[�����UsN��|��㔕���kcn Q�H�!���荇�#C�IY
�n'h6����E���{&bc ʭZk��*$�:fDE_a?-����s܂�� O_=S�P �lt�xp5֢G�� �̹~_��2HA"4�ms=	��^4E������1�(ֽ�״��4��?�5�]��T�S���8q���]��� �y<ֿF_߱���*�9(��4���D&�����P�xs\��E���|��Zb���_&���MȪzk���l@-�k<d�����a8�0����,�� oWX_=��ZƵ�Vѐ�s�ͿH�WD \���ػ�Z�Ǖ�I�'�_��V�D��"<� �Riw2KTi"хR�>�i��PI����gS�����`~��+א��.�ǲ��D��δ�͒3}��2z��K�B[�zjz*7��Υrb�N�،�,0���W�����M�:hA�Ỡ*{�����mzޮ�jH�3�	['�@�.}��sі.��S}�V'�/��>�s
{�)�I�v��q���bv���_��"���4�fw6�l�4{7ඳ����<^	.	F�~�ܴ�;��S$א���<4���c�����i���rr~���;�M��5�e�r��Ñ�����E�x]��׃nǶ�1�q2x#F���/��?�]�a�����M��۟�;nIF�~h�{ށՌ+$��.�	b�SuX-�l�e�avZB���5�oH.�2���)h��H� |G��I37�F�W�n����5�Z5�DN�9��[N�a�2��Re�� B�z��Rqz��ig ɘ�N�j��f����o�:m�1��]FW�Z	�3�D�ܘ�O���t�}BH�ȱ7��Ӡ�J�9fX4�x~�Rg;�wj6�H��t�(��n�mvՈ}�+{~��D�'�v�P-	<������B�˺8ͽ��6\���5�#�{M�0K@"Qǻ��*�U��|�����r�u&	��V"���=r{�h�d����*�@�J�����9�I�-),o
z�����R�M��]�K,����FJNi��y�%Gk�.VQ+�?�12f������.El��O��������(�����/b�j�2xw��m�_0i
�_�\*��7FEC��b���g�m��[���X�R�/$��<}�9!�ƭ����%�m��:���2}��_~{B~�S��e�p�䭙^-��N_�@���0�}`�r��M�	��Gm&���A!��� �W�ZnK�æ��zݹE(������qm��647;9��C���c��8R��L�ƺ�l�d
��I����X"�@o	E��c�pJ�E!U�
�c{�ѵ��K�֍��޺�Ț���3:��e���nOC��KO��W��G����5�e�6�
9�{��sa�P	���?Qݩo�.��+	�=������^[�/��rҖ���[>���@�i����Vu95�>���U��$���D�
V�4{��ј�$��B)��д����`��j#�΅c�z{�^k�b��O�(��;_ZȓjA����c�1�w�|UceF�����³�"�p�8E��r�N�VB�=��+�t��}����M��<s��t����iI�a�AX´{y�}K�+Z�o�cĂ���t�v��?dC(Ć�=�o�B�-��L(Ftw�SwnR�P�'E�j?�:�[�-���HE1�����y�fei*�$��<�r��B5p� �?�4�M��=-�[�%Lr�賁� y�=�V˟���ӝ��J/������ITA�߁p�v(���������ɶ��9��6�VCxS��	��w�=Y���]K���X�D=$(|�q���(��"	s�lI9���E\�^�M21l�2e�%�r�I̾�ŗc*�)�����Fp~�r*��C���lȢ��c�C�3S?b�&��z�w�I�T�X��-�j��8�mヅ��7�X�. �:�h���.��5��.k�05�ħE�o�v�$|&�y��T"9
5�ߢ�}�t�$���E+��;��"�>ɇ�'m����80-���	ґ�O�Dc��Ž�ܿsǇ�rXaSh��:�_\%��,U|�L�r.#@B�OVT+����ؘ���'�V�2��<�2���o�Bll��B$��@�0�؄~�f�
��w�����d���ł[�*4i��-��8cX�;r�jӳ�� Q�Vه����Ѳ���`b�M��g^dܚ�J^�҃)����z#�[��p��i))^,���z��b�<��i�?�o�@�&_���r���SUR�� 5�d:w.E(7�~^GՀ��	09�N��iB��]n_��j~�z3��+������[��͙D������=�r\un�����zz��L6M�Y5K�A�|�&����N�v;ԙz{,Lb��A�</	�/�x�e�/�5��ݽr&�Ip��Л��䖽im�Z"����?|d��h��Mrҙ�	0B�ǲ�v���l�cCMe������VP��$�P�Y!-f��.���,��.�Cc*�VX�������O��!&�:�Ȉ�v����3����*#h`������h|o�f؆��dZ_�I��@o4��W�$��H�+�4̈l�Q=��R�l$j,д%^���)h8&̯��<37��Xvt�5����qѳ�&x�F���'���d����5ْ�k���E�6���EFk�#�2�~�S`�[����w��'g�N'U3
>nV����^ܪ���Q(uU.U�h9�}�&́��]���GTȞ���1>����)Ž�-0�]�+��O�Q�Έ^mjrW�x��������|���G�もS�7�r��\�R=)z���et�x�ld�D�T�t�tl���d��7<BI��� w.$ItP�2��7�:p������ּh���p�h�{�|>����A$��{=�U�rf|���FЈ�逭C\%����E�j�#h5� ���W�;�ٯ�w�;'�=�V���)j��0-5l9aeG��[h�)�jd��L�����ˍ��HQ�pO��������:(F��LA�>��-�ʷ�����Sx�f�Ԑ��`a�
�&��ϟ#�G��BG_]9/��12�e�ӑ�g� �C��j�rH�M��j�6A��5=�ޗ�~蓘�,)Է�<׺χ۬�ВA�:�h��.�c�νfs�WTQ���pg$����uVK6�4��F��&B����ϰ%���"��?M�2t��]\�
0Xw��N���Mx��Q��X�$r�d=��ޚC�P�Y�r�=��3�����&�2�\�s-ϮN��j��uvX�p����_~�H ��[ο�]�&�uSh7�pE+"�� �o���Ѧy�Wʈ�k����"�R}�sڻ%��dQ�ʅL-�\M��چ���1�PH� w�����4����%@^]�N.�y�$�2s,$G�*�DE�&x{F���k��Hޒ���[&2GKZ?4�yh�)��&��j���k�b�~r�=��+U��׆�(�՗g�K�`w�6���y�f g��R�>�3�ns�9ב����i���~�`�A�l��I�.A�ME�k�����Qt��/�1��h�� <�e?�V��@k#,)E.���c�T9��P���L�{�@�&�'��yGPD�YF�P" ��m��ZQ֜�l��+�X�tyS7f���� Tl���9�m{�|0�����ܗ��>Ԃm�6�1"m��_Ƽ�z����:;|p����{Nɻ>�h)�w��t����OGdr�ֿ<��ݿ,i؝R,�~��$ӧE�u-�j��B~�1>��ZElG̔>%���_�"8ر#1W�)��|��ߤ~�Tt~8Q��4�x�}R��Z.!o%.�	�v��˱6T.������¶��8B�| T �)AZ��$�{�Jt��h���#iQ��,b�Z�%�ϓ0�O�k$���F����3�]	�GC=�̏��v��=P�ӯ�X(d�Tis�Y�j�1P�L������[���C#?$N�PH{��H��x뚿��C�$�M�~���el60pG�ί�u����3��x�.��ն�izy	�j��ZE��Yم��!>��{��N���S��r��b^�&*@�&v�\�63¡�?}�������/]|N����}����Lx3��z�T�פU~� �ό��:��)��<��R��.1��[�����a	�#�C�Tf�����+�+��~dp&�����?-`	��6�}=�|�?�)����E�#�L���X0��.�g\jTȶ+��X���g���[�&㨱e�ҟ��d��u�̥Lod
1=%Z���;���w��2�X��H�D��?L�S[�C�Y�(��ʪ�L��œVV�gw f(�F!Mk��|w�*\�)�ߵ"'���t%n
?�Ը��]�����5�*_�
����#����̨�2��#��`���H֌Kњ���Gic��$c�M��x*��/���+��/$�	�T�_ ��ƪ�[!�H�b�KQ��vچ��g}Ch.�x��~��.���0�5J2�JH#����p��l�i淙|�ˈO�tV8������Ȓ=�����=T���������Vo��0b1Q�dg �N�zͽ��&���O�0}$�a�t�Q�c	�ůᐬ�����F�Ȣ�6��'�#�:"�Xld.@_��J�V����kf��u����h(f�){~ <	��nH �푻�#�C<Y�~><��r���k���c��H^�5{���}BG����H�g
�!�;>�~�p�.�3���g�O&�#�/��d��W���G�dc���PLu�Q���1���f����fJ�����ut�GYd��i�6rM�C4�F�w�DJ��&U�tӼ-��u��1��@�1�I�G>@��[���S�_�
�����0�����N$c��9�˔xƨUE��oBZ1�-�:��]��+��n�Q��2�wU�^�
?1�Q�F;S��m ��g[�8��*Zf��a��ۺخ�����:�u!��,��P�Xk"c�T���e�V���*R�Q�J�GX����5�¤��/���Q�c�4���g��6�?~Ǵ�q�J���גK����'�Z��b{���uh�"F!�Z�lH�/%����ptQ:A��lL�y,�<Y40��eL+�E�Н"�V�����W�fn˧CLT�n`�5���'I�z�F߅���Ţ2�b���.�@B�ó��@e�p�r�Ҏ�nހs�*?i��qags�^O$�;i��S+��p25����b�$Ih.���e������]V=����9�A:)�4��pS�KqQ�l+�~�1���a�9�=:�1�~} �1����a�ni=�֢����@�	g:I6Zf(O�����)�4���Ŝ���!���Sh!@^tܯ�FK�W��������o�i����Vw�9��x6G�wE?
�^�B$�y��}v�w��"�W �"�&�Z���;R0��d�����������eC��\S�?�i"��&w���R&�@�|��WCH����xvu��u9�V؊�"����C����Y�����_�V`��z�`�O��V��wyR����׃m��w O�௜����zJ.(P�W�P���wB�ŻZ�SV�Zw^H�~IBi�ɺ���.�Đ�T&`���Y��YC}�)��h��}c�8������n�K�� Nj���IMK���t�jg��!�u`j�D���n����EM%<�y�7J��4��x3���1O�[�����������o���ܝ��1����Q�xV��ēNt�$��]����Sp�|P�Lp<>��R��~ap�1q��
d�|q��v4h*a�Q�(f��4�ِ3I3g� �Z�+�Ǯַ�=�g?6e�w4�����H��L|e�	����q�´A�U�H�+?r7�,���όhD�A5��q�wM��yNLǷUA��TO�
Ӫ�#�^�r�0�:Zq��K��rG=��VG��p7��z��N_JX���5�+8�GV<|ƌ@��?s��05i�p��x�+�3�^����N���f�Ru���b��ؘ�^L�NMU?��=�ӕQ � ����/��N1GL!�����L$QU�� mĶ�;���JW� ����M�y�&ۃ�q���Asv�l~��9?Y�s�?�&�K���H
�d5*��o��������7�ͬ�uc	)ia�$�Uٲ�f{oӺ�:6�.��ϕ��5���Y� �m���U]�`��P�����ij����2��n�k�Pwߜ�iQ��=��⢹{[����c.-&=b�|�)JuC��ګ#Z��֬Sʹ���^�-�����n�Z�vM�';�w5V�����d���S!ų��2��
B���o4Ϧ8���[, ��tC�B/�E��0�S�3��	�/(Þ譴N�Wp�HG���/\�]�N�V/bQ��K�V̝�(#+�`��s�|��E�C��u��G�9��.Q��>J�_5�:�hH��4�2�-��{)Q< ���>/	D!�h��G�* �9��I��@n�|zSn���g@
�}��ۍ>��h���*��3��C�����~�TVb�zgH+�N�w w	�Y}����xU�!��A[y>� LdJ��nW'���w�1%����Vy�5�7"�,|�c����1~�GX.�8��ܻ�����5��QC`i���V�#��fa�>[4���g!${���7�`B���zMTO�A@�^^��-�#SN&.���Ͼ��B7�{-�%�j�~�ǎc�'*[۵��Mˌ�e�D-�ߚ�SYP)C��40
ad]�%y� $��J���B+_x��Կ�~�|�}��H��z���>����mȆ=��j�B;�g}K����`�|�e�28Х�ZvsXs>?�g_9R�j�AQ�#'�[7&�i�]��,v�i�/�UP�{Tх�����ѯ���k�Y�g�Z����i,�+	��A�����#�0�?�L�m���$Gnn��z�����c�-�#|��������f��#}�F�Wy�[�[G��5n��*L�H�@ n��ϓ��w����:p0�`d�`[�=�w�3�ãa�&�F�l���\���l����,��~qE+���2�J���<]!ʭ�*�g�h�v"V���
=��L3��a�Gxo	�(��iL`Ο�H[f�;����pr��m�sB�` �b&�\�u #iGH�����[��=_ɩ�!�� �+���,k����'<��Oy���H{$����r Y�hk�1�dY�� j��_�XBJS�e�V
8�2	{�8���3t,���v�lp0	Ҫ�(嗖����i�,�H�!���]U�{����Cʱ`O���Lp����=�b|�G�C�6�7�{H5��4�n�p�J���˪�[*��՛���j4��V����2�Kw�~d�C����iH��ZW�3?�i?-	̱]݄��'\۞_l��X;y�]�!�A�U��� ���h�� ���p0�/�&�ِ�k&�ߛ����Su6��U��+(߮_:�"�U�b'��5�a�1��W�!G�%�Z;��i���3ow)�f-���m��@���ڇ
����	ￓ��ɿ��r�d��l��C�œ�('jQ8�e$O�z�����W�T?z�d$�X$N�f�\�`e�ք�)ț+�����P�G��`O�-*�b"��4X���כ�g�p�)�'07�T��K�$�zYt�&�;�X��C��L��*��Y�� U���fi�A~�G9K����<'6�D�j���_	��"��5�����x���]%$ ���F�&g��6k���-���Yv����]�G�#���	�H_nX�w���&�m2+�" s����Ջ�������8�/̻�����S���U����64�#�B��ʁ�ݤ?�uLN��GW,�DNuI�":mw��Nzٟ�yK�ts���1i��i���L�[a=!�48��l~��&�ZI.$o0�7�D�I\.`Rֱ��j��� 黯e��_I� �v�6����I��KI+��v45b_@/�_dw���]��q����S�����Zzڀ����Fj��3���(n������C��пY��E-��/������ss�'d��;p]��d�A���˯���j"�x�i̫�"]�)��fG�[i�P�DިJ�;�T��h�糂x�=�̜���?�4��&'Ġ/O���ǃSѡ����)��=[pJ{��� �w2ˏf�ZTTU��Zf�K�͓Im��n�`��n�[�\���4-�?PnȂ�y�;Ի�c5~�^"_v�%��#�K� ��?Ji"[��Wb��_w�� þj��Tʪ���1*�M�s\Ɂ�y��`�Fe�8��N^m�^C�� �*�'�	���
�)��5��NP��E��`s���\[O�(%'�Q@O"u�ܖ��+A���E��e��hJ-�c�.k�.-�дnh��|����x�z1>������(DpQCt�Q�,��V����{`e{�.�3ū�z"`W4�E�>k����%8O�cb��}���/CvLqg��P�.&{�x|�����k����O��Z�i��3BF��27~9���L,��'�i�tJ�����}�h��>�ES���`�($OCi:��f>��}�hێ{
_z`V����J6!<􌶽�ZJ��_�DUw��KM�����A��Iڨ��DHJ�ڭ�V/_6IV�K���A�sz�˘y�JJ��UA��E�9�&s�@�F��N��1xD�!�bwyU�pV��x ���(	Ȩs�G��@Z�d���
;|%9�\G�c���t!�U�Q1%��j[����qS�i������?��8H�^���֮�Cd������q�2���֞�D�T8ӑV!�9?�vk�-B�m�w��Z8�Q4����E vKq�p}�z��"����r�޺@�٧.��i�v;#�E�J���h��V��7�Y%�w�gg��&��v��t��G�<�rK��y�|zL
d����<��(�&�V��g�˓�5�NųЫ��L�6x��%g�����>gz���� z�WCoq/K*�����~jq�a��4�~޹B���'����?���N+�Θ�qBnQ�B�G=��$�.���K����G��C��ւn=�#�7��X�c����@L�$$���Zhſ�!�1O�;n����aDF+��!��������tdv�o���gJC]�����H���a`�l �Wn�1k������#�C[5�/���೙	��I�v-�VcNPPj�*\���<��{G�����]� �z[����J��K�!f�R(|���0,���^�Xg�xtQC�\�=�S��J�i�ql"�*rWL�1;���+��k�
�S�~��qA��7@��e]qr�mzg���Qr���õe�W!�ޡQ�g�Z�� �G��_��/���y���Nw�.��"~� �IY�y�EA���$b1ƙ�8V�P˿�y�d�{d�λG�!>��u�`��itLJٹ9➅C��4@�v� �
7����슖�`�ai=��9�
�n�4�n�q��rt�G�ׄ\����VU"��(�Y
�f��q��n���N6}�G׵����/N{�#c�U�L��t��e�)�fy4r��j)�>ce��BRPg>d���c=�$a������ڣ�hc��{���)��&�s!�n�
;k�^,s
�\F��!�$.��X�_��Ú��p�j�\	
 \BD��K��]G�0A	j��J����G���Jy��o���M��j[�!���ͺ�>U[�G�����p�U��Iq�Y������q:�SFC4埓j|�4�5��vp�Ŕ�38�zC���-m*�G��z3����fh���S��R������h\B:������}��!fj@ST�z)��3�S)�r:�C��d��e@q�c��5���hi^H����iݜ���V��s��of7#s�Ά�3��Own)_�YI ֖��oa���O�!)P�&^���L�V��lL�2�ôט�O���2J��^�z&Xo��(�b�\�
	�oB+�74��p��z�rs�᫾�I:��-�JH�k)MRX"��-;��f����O,IGO&.��W���Vm'�^'�G4?'�'����@���Ж9e�*���S��,_r<5�t�3������c&{*UG�ԡ :HB�_u�Ғ촵��̂�SD��p��o�]�y?��%Z?�F�J'iu7ܜX�-��
D�t��řA�*|J8L�Rzŧ[R��{a�&g��Qx�|����-����ǫ�;y��Y����5 ���`6��*A|t�?<�E�y�zQ�֎�?��?����f�c�	���'C3���N���=�,Yg�f#�Pjp�H�1�AS\Ȣ���h>;� d_w ��=?�����u�T�r��jV<�p�Z޴�-?E8miy�?<�@���%|i�g��f���x���� O���D֝��EG�x(Ɣ�؟O{P\��H?E���$��ؑU��@g��ֈ$��;Eb Kb;�@���̖FD����yM�v*$p��%2�\T����㊛�<To���@�E��_��h�V{D^RL�(F�1Z�8��+��9֎�*�g&��R.y��˗�h���F���æ�4�Gj�we��ûVl0Z�"��I(�R�N�Wa�K�>�;��6²������� q�� ���m���]����:�j�o@�r����|�<T������ ���b@C\zㆈ��K�$3��<���9��Ý�YI�����
�`���Q��sȧ�ρ� ��H 4����8��Lz�fO�[f��AV�e��t�^���R�?Y�����Bs��(�t���m����֚o�gp�㌻i�3乁r�������]���20+�-�B���/yw�%��l���s�%�8n.R6�`�b9C�s*��..�rO�tM͡?�9��i�A��?�F�� `��SA�Y�>)�	Z�4�Q���6)e8�Ҧ~��=yOʺs�D����7F4"e)�"�	9B�w�6�R����S<d��!��Wg��0������W�e�T�*V���Bl���ơ�f��g����ww�U�����Y�)���.S�/�,���b�9;*|E0h3�,��k��{���U^]D2��܀(P�8�gc���5�O�.g5<$�Q�sH��Di����*�!�Ž��$�?S�Ϡ{k����w���-�K�^T%U'K��lH�zd�[
d��|�ogF4C�����Mh��G3)m�����M�"���y&Ny��ڽwx*��I���@���
��=��0�:W�z��)�� �NB�b�O��1�q�q��c��}�kӒ
����~���W�1���ұ�-pN��$XTD�8�@Q�����E�AAu�i��P�(��Erb#ĳ`��QS�DAн��y^˝:'�xj���H�M������rӈJM?�~�Z�E�v��4S�,9H[��]�P���j LWIEw����/��4��'n�p[AWI�I�e�\v��>��E�ŋ�S��T�K�f�婠x�[p�hւ�a���"
U�a5xʓ9� �T%��<�n��	
{T籒X���򇇽x�Z�e��dRZ��3%�>���r�.nM��t7̲|�q� �U�Bmz/wBõ��̺�:�z�^�9��=XZx���V�cN�0�T��Y������ ������m�02�T�e��7��}��"h	�0c)�'���c��}�h����;�����8K���:�j.l�34�VTqQ�� ����Z��d}R�M�R��w�ΔI��%�El���C�Y�O@(��c�����)Y|����dKctNϲ�~��U�xT��=O�5R�d�z���Gp�"�9g��%�L,�BskV�ꊲ��I��)��L�(	Io\�W�������G_J ��W�b�91�R��[��I��R�tߠ���	�A�y4��A��_6��W�5�FM E�X=$�^y8�I����Tp��H��^��]e�Ǖ��t�[B-��E�1Y]#�c���s�	�1�)�ˌ��n��З��Z,�	O����r�Υ��"�s�i�3ĳ�M58�֏�5	�A�*MA�>j\���ϔֲ�O�E�U�0ˡ!ʩ��|�R�;��>h�
��J@b�J���@�IA1q&Ê�3!tff�v!���������ʀ�,;�$D���`iC�Z��<���x�Cge�%���r�"!r��bb{*P^�
d��	��)��������5hLE���jХ�/����}���%N=*U��B�F/��u���5d�`5(��&4����+ԋM�~Oh��;�� ��d�Kw�I�ы ��O���]C}��,~��g���pZ�����,?> ˌ��|M7`�S�f�=V���
��Hv'�R1�Z--uy���Y�I3d�8W3�h�Sx'.l�J��$K�։����,|��G�H_�������n@>ê�hM�����F�^ȡ��
�t|�t2�z牦��J�����]w�TE�[DO��I��|�X_<��e�S8wt� ���M����`�BO�-A��n��m�ul�QQ���A���No���נ�`���� �g�����
��h�J��Sϰc�p%i,�>3����gIGT��у-1`(��X��]�!��7�w�Y[$٬�a�0�~�.i�[ϏA�f��cNE�=�^�I4���v9�6�~zU
*{p	�0��M`a�[IR�Y��-�zC��J�(S��M��W�3��D#�Kq��U��:�,�4tp|v	A�8s�f�R�Oc�m��8��y�R����Z\�K �c!i�?��xݑ�/�b�#h�X�!�@�D�T�s�g.���uM�RR�sq��
1�CJF����w�-�u��įx�	6Q���%d��Urr6�a�W�x�c���U�_ȕ�u�EU�#��z�q=Ɠ�)�"�d���!���c�������R\��o��dᾑ{&!jW} ~�[�j3J�QX�Ҳ7�Sa]Q�{���㯂���^�Kv}��� %����i|L�.}�:k,UBI&��d�RO?OF(��5����MD�&��@���ڠK���i��!u�/�s��F�}� �߸�j`��y(�����%^�X�Җ���?S�c�֡���VQ�Œ|�%u�s��	��cgG�tm�����$�>J�p��{o=�<M"���d�c���ŝJ=��^0>���@-*d��X(��jC��i]���?���&�g�i���E>�3y�J�
*A#vA/�ӥ���љR,�-�������&N���Bg�	�.h���L����/�?*�w����	���UF,�3s�_�����yrd2��� �E¢�� �Q}Ea��GQ��l$i��I�1�9�es�!8/3GJ�bC�@f��]���BM2���}d�
�bD�;4Y aE��)�����&�79�^���f}6࿫��P�D	�1"���fNi6���p~�}���8�U�.���_�J��w������Eh��hQZ�g���dd�̭!r�cz�vn�1?�)u��(P�2��7g'K�Vu�}�F�Q���lJy#Ӹ�M��Jv<0���Z��ѧ�x�~L��N(}���A���ٕ��������ܔ���"-!��?D}����:DZ�}mg~��̇�R,�P��B�s�'t.����$���UX�u��N��r��}��:_����g>��$v\<�d/GnQ�|�x#R@{(�|�-ܾFē6ݲ���C-�)6�	#a�S�6W90�:�S�������G������\�M�R؅��C��U��o(��i����-�Jo%u*�Z��ƣd^���>���t4W�7&�g(�1m���Q������R�*�6��XE��l��?���Ij3�"k�T`jz�Z<�I��W�Z��$���!��U��Ǣ�_bH'�<f�mD�*�7��X:��/4��^���>p���4l��-�e{�`�̃-�T�����5���B�hE��
{,� Ct՘���4���j�Cԏ���9��g ���@șx�?�Le�­=E�x���J�D�&:���3�S~M�ef]��<���^����֝:��u��Ce���!:��;�@4x�f�ϡ��J'f���d�;�F�O���7P3���o�ݕ3&�=8��}�t�R��������B��E��p0�:C��{�%wl����@�H޸iQ$�½���}�t���k�������k���t9��wD0������ڨj�9�z�d�QUBrp|1_Ap��.eW��n�~�M.t���WT��\"�9)��}�_����灠�m_9�������)-*k:�W[z�+�;�#=���V"�,BMy�K�\X9k��nՖ�+)������.Y,�,݌�`Kl��uy��C.��Eˌ0���D�D��pV�_�}%���#����uS5�'��_�g�9:��%��D+kJFkR`~%R�/�P������xȾ��T1���"E�6L��VǸ�DC�Kk.vh�v��=�d�2)]�=�_�9�H ������v�j����5h�˫(KP��4��B�W�Z�7�0i����;�ؠh18�v����QF�����׋������%y�z�m_�R&��mq[T���_�|l_���Y���Ze �ń}l�
5�_���W����pg��Up, s�ct����n�H/*��E�o���>�����ʗ/Z|,^�Ej߯D����M�DBP�cWT@�{�%o�.v�5��Q�
���#�.Z�5���:��X49� q��t��r3�Kq���O 0,t4j����t{޿@�U�����7�[��L���,$;�Ij��r�[�@t��l�Jd}Y���zqE�M��*���ސ��ۢ���F1@6]��&�Ɲϭ��O��6�t�'F�0��E6'kd��ϏBW�����Ԁ���gޠ6�#�Ԅ�|380,�{�Jw_�ZQ` o�l������Y���fiV��L5�|������W�$�{L*c-c�5`��~0��[6��������M2�O��#�&�Go��]���;<����c�';y�Ыg$p�eޞD�U��JT�	O�`�ל}K��^�� n�f=9��鵘T��D�3�%\E�ҏ�Y��U��P8�c\�$d�����I�n�଱ӡ�Pi�)��Я����I��/u�h���b�	����]Á׎�b�m��$i�̕'I��b��F�ຎ���D�aSbbuD��:� �2
�W<�H��i�l���@T�>o^"@�?��ōi٨_H�	L��ך#�7Vk��x��eo  ����
K�R}ս��}_��b;vif��}��n��2�=��:WD���s����Aw]�1�H9;0l��;��r���z�A�1m�熹��"s���m>�a�k���S{[�)<ab�~�f�0F[�Ӕ�,1�K7�UBOhL�]��T�"�[��+��5���hP	�p2jΛ�ɓ۠f.N ��V�p	����Q�Z,�\˕�����n1+��.QtQ�UvvS�ՇLy��%ʥ�J���M��&?�j���|��m����7���x���]���I�V�2($��#�#(@Oi�";W�_j�i�?�A���:�*�]j0���i[
�	�f\H�<hgAO���a����m[�%%]̬�D@H���d4�9����	�@Wv#� �{yB�U����Ӫ?i��G#}���MZ|�H�.8x3~�	�Z����z�����e���
�Gڱ$���}�����ܸ��{1 _>c��<��H�Pc�X�5r���)�����Y(g���ֿF>83����kU"�N���\���:�؀��#w�ؒ/�b�%f˗�y~�S3�v]/%�HԱOe�H�kI���F�jj��u��\ ��(9�ǡ7�}��N�����l�	��9k�A��Z#%b����h���p����ǇR��j.\i"�z8��m+�k^L)�]JdhI��+�O��@]�%`A"&d]l����}?�Co�6"���ԡ�)�˜���wĦ���sc���U�R��AK[%�{��y�:3Ƞ¬��#
��DIz%T��<��AL�N�lr�i�j:!�CR��@	��
q�n�Aʱ���i�t�@F�w��:{c�{����U�,	�&�����> ���Z����9p�5c����v��l\��Ij�\se��H f�W� "N��{�-R��`�[+��":��6H�&.���!'��X�J�;���-zo�p�A�������MM���AȥV�� �S<�����i�<����{�QS��}����ը�Ё抒�b�#�Pl��6p�s5��~]'>\6h��wP��������Յ�T�X��G��^d��s,T�h�O7�%³V�E����3�,��x�}D��VM-?��"m�)�o�Q�u�H��]q��m�� ��k������j������-�p1p���OG^]V\E��.�Q��iܗ���c����� 7� ��������qb�C὞ȵ�QAw�ϔ[&Ͷ�߱�j�Pݵ�~�vɒ�c&a��Z"���}2vr_5��EA���2�_�c�HC(�˝힪vQp�[��ˤM���w�����a�(d��bXj���?�AC��ʬe4p��,�J��ſ�i�]ה��#�t)5dfM��5U����Ⱥ1(�F�S��Ϩ�"|�4?ӌ \��f�MJ۪�	�ynL�\�<�4a0ߊ�X^y��3xy/�;�Ԛ6�ъ��h�]Ѳ^��a�dn��܊��\�Cb�z��{������[���HHGd�L�:��/�MD���kG�x��n\����1�Ȼ��=�X����GE�y��1z����6��T�â��Kͻ�"dt:�l�����N/B�c�\m�j�H�AD��׏J��BL��_��`r����ql��[�ã��#�WT�0�G�{^��_�0�%��������a]�dզ�<a�~�����^�c*GHp1a<ځ<a��8��M��	��y;��a�a
�0
a'��N
Cz�%����m�]��D�^S��*d�q�a6�n�k�b����ak�.}���D��>��j�0A(�C�JT��������<���ӘP���ւ�-�K
�_W��1���ﾉG
�S�m`�W�y�_�лH�*�_�����r)p�l.�/Ʃ�I�	�L�\��V�#�Ͳ�����R��Q�Q����ڶߚs
lul|�5jp��9y��HW��x�ֵA6�E��	\��+�����N����Э�g$#�Z�u�ˮ��Q�����U�ut8����~jn:������y�{XWyj˶D�Z
c�R�0��q��Љ"G�l��F&�@��۟<r��I�40��8��0�}��1�B�TQ�QJ�6ƹ���cC��m]�?˟���lJ@������n�kz�]vbP�吡Ԏ��ƔQ?I3��t��|��Q� ����ܬ���pi�11q��#p�"�*J]$V�!�Z=q�o��e��g[���޶�t|D�^r峳���9�~�,n+n}��ա�Ve�a�g�ڥ���(�7r�2�X�\x�!� �+��ф4O���Iꉾ�M�R��~ ��x�kѫC��y���.� �!������v5��;�t�N�3�m[�g��s%dj����gۭ�ܗ�v��5�Ӆ��44B�������~}S1�2�A�vm�~_�BR"�������b�,���+gN~줉$.��L�2_���򲏁�ؘ<r
�h*����b
{���p(��M&���;Ħ5��i�'*ٹZ~���Cҷ�KW��v�'6:>�m#�̷O� ��c&��l���G��˥t��`&sNǘ�uqf�S��x�Z�2�ƯRd��m�n@. z8����H��au.��ϱ�I�}�"�t���Hg����18�q˅yu7��&��S��:�]��[h�Ź�vر��3�N��'f�ǵ�ho���F�l�y�D�Do(YB�U!Bw�h�oFy�����>jMl:����#ɹX�l����<K��fΞc_Pz���%���l�ˍ���	O2L�.�ҭ�%�Yk��z�y�P�YF��o�p���i_K�nL�7�mr�2�;LG�&����!@�JW�jM�YF��_��}g�_�j��0�j��t�_��
�4�tt��zf�VŎ�K��)�W���n�O	�Mr&JD��9�$��,�lZv�������(ױ�O��b5� ���}�h�@ώD� WZew"�����I��!ʶ����R~%���?�4ek-�L�&py� ��0�J��a���9m��F�^���9}�N�y�M����Q��8 +�]¿6���M�БH�Z�8�{��,:7\BR�ψ��x"�6��`Ԣ8�ݲ�9����N��1MՀ읭� ��Tg_(?���<�.�� �����c����A���hxjt�/I�Y�(X+�d��+u�N�
�'�)35g#@e^��2K��+����)r ����k���Y=}�G���P����#��a���;Q��N��@=[���S/[FmlZ���)��æ�0\~7��"I^���8Z�.��"����-��p(z� l��_	���� .���]��ɒ9�n@�L.��ƀ�ɛBqԟ�҆T*ro�B����q�~wg�ЫE8>��$q�I�ы���CJK��}�H�Gi��n�<r���Ň��t��8�E!��
}��Nn��ZȺ!�	py(|�(R��B?f����$�,7VF���ľ���_����'r��;_K�"��웛J�X�OQ���v����Jb��Պ\t���*�p�@�t���;�t����i�*�G~!�#Ep�TγEƞ�<6���ML҃?y��'���~�����X*�����?deL`f=�G�Ô�x�-�`�Ə��y.�����#b쮭�Ɯ�3K��R�r�bqGM���n��������9B��s�\]��B(<��B��U�nU�}�8��!�+�N?�B��+1���
!�^�8��%�i�W_(þ0����ђ�;2nr�����X	D{*�u���,�>�r� �b D�cp�Ak�j����z��6����w�n��Yz�H�%�q$i��r�t�w�ue,�K2�����a�{!F�ښ9�"��䎼1��wS���R�r�cm����y�)�c��$yF��%֩ N1�e*��O���PT�\�Hx,Ǐ�E8��L�o�3�|�R���,#0}pgf�*��M�o{l�8�#>�ӆ�P*�Ǎ�6B</kGHʺD�;%T���^yg������Sg*��k����C� *bːß8�?2I��m�NN55A 
 �1� %c��W˰���|�	�vA�xS�nr4����9N>p�1�#�;9��o����q5S�5DJ�xhm�#x*�Tlh��3�ֳ���f��A������&J,�5)��q���G���mђ�!�ed��R0���O�����E�Y�f���G!3�>�C2�S*0�U/e�k��|b��-��e�h4l��A�>s �.m�6�/*@�ݺ�jttc����]N�,��򬉬y�����b����Y��B���B�8��[��Y`�ɺ:�W&�[>�!m���0�RdG��/�]~�����$I��=��GU>�bN�B����6�G(f�Q��(�<�J���|����PN?Z�q�Pn���#8��/�`k�Tk��3�V���f�ط*6Z	ս<d��6>��2QX��k�ԁ�3��2�J�J8g=Nt�.�Y�����aA�D�,/ؿy�B�U�9�͎B�i;��k|9��nU%��'�{�ܟ��c�d���ㄥ��3�H�g<��2�Μ�����~w��d`�̇�Y')?����5��-L���D5]�z���_����� 1xݵ�&�Tṏ��t�_�ڣ晲,��ʟ��+/ᰃn�)O(���|���O�Sm0@g�ׯ]��j7|��3�U���V��Y���:Q��"b,����\|��W������/b�2:Y()�v[Ho���y�ᦵ[Q�+�"/r��s��P��cP-�:����>`�����b�x��<��.
�a��<U�c%��H�j��wﾆ��>hp3������=�+���s�͜k[S�V/�e|���?� FKY�$u(D��4��_��K�o또^�����Mw�Gv0؜ú����h��4`Z�'�Z��y��.l�,��e�̃�v�Y���N�.�b�f����z'���x��A;N��C�ȋ�Y��ަ�f�'�]�ߐ"ov���_���,�k�T���9C]g��j}��V�`��!aw�� �Nd�����Q�JJk���A{nu���M�y(�'�,?/� �.!�?�F��b�Up�t�D02�5S#�|��=Ҕ'���jB�Wȡ��?�bI(�bx8(W���Hg�W�U?�V[Ⱥ�(M]:�!��-���*b��Lx1ȏg ����43��D��6{�^�9���~M�3�~�4��&����O�h���{���Ǝ�cU�F~'�=�Nx
���{�w�ÓPJ��vV���sνkRޓ�@�GHݎs;R�H~�lqm�M��d�p>�F=B�n�I�Pn^Z
A�;�R)%�ɰ�ᩜ�*�$��'�}ɏ�CxF9�o5�e��n�:d��r�Bo%h�e���v�K�O����vo��N��q��3<%���x�@x��!6�&������C�e�(�7m3�1L������C��ߕ\��P_��/�N�	�%����aσc��2��L#����^��Tg��.�H��a�D�h�G_�Yz9<�NEb⅙E2'䄀��Q/��d� �߻jK����l5�琖��-�9����{��/,w�Ày2���
&��x��r��Vs�V`��$^q
O�0�w�?��e{��Z8g���J�m� ����Y0p�;����)�*o���N��9���i�}o�q2x��P���������"�?���Ԥqo1wp�*�r�oFw}�����E��]�j�4zUuj�a���A8���w�������Bl����}�����m�a�����s���� |K	�cGe�Χ	׌]y�K#w$'�� {ÜҦ���b��]�� �Lb�D�X�e�UC�T,W}�H�᪢iο��Z�MAdp���Զ� 1�3�y�KW=��ÁWr]�<�F�EH����pǷe }�}�f�a?RD�i�;}Q�F6Tɸ!��5[l�%�2�G��i���~ ��&f�bX�g���(�eb J��Ӳ~y�1sm�A}��x��U�I��Zk�����/�/��ug<�m?��{A!�Q˝�nZ�<IЉo����q�zem�D������ű�����V$�+�Qq�6��HL>����*_�ӎ�Єg�1̂��F�5j���9���q�����w��������#d����Q[!`���Hg5�[ū�>2��E(���{��i��yl7�`RS�a+{�G����'+W�l��f�p�m/�6��&�Y�zz�:�1`^�;E���O�ǟ��<�΃4�� ;�R��V�z2`�h�Q|��/������l@���@�J��)� U�s�=�� ,�/�P4���&�-g�!��2>vҘ�p�5�9�DQNr|g)��X�l'$-B��.����j�����ؙS�C�ko��9S|�T���ms��&n /g�Z���"�}��Rf$�䫀�Ȅ�f7�~�o��|S�0	jnZq��S�6�џ���3���ǿ��BǇ�[����.89�'�˔D~���`�^xT��@O�5\04���+�\�6>Ryz��8b^M� �y��Qr'C�7���׍�;yŞn2Q3<���m굲�E����^m�h:�����IȻX)�<�U�C!d�����f9)���gS�4@�u4�������g���(F����kͶ�}��[�~T�[:�j�ü�)�`�������������  럘�sx_87V�j���T�"t�^�,"�*���XFѱˎ��BnÌ��2��r<ײO���|.�?��=��C+>���C|�.�2�D�����ry'Oݪ�ȉ8���M�i�����	����@=��H��
̹ɭ��5�zǯ�o�Nu v~�WJ&p��.q��[ٛh���
�N�Y��0�¡�0d����f4�V���F$	#���#]?VZ�u�c�!����{�b�%��������"�&�8�Vu1-.��L'_��~R^WOO=���B��}:V�Lu��p���m��vX@�˄@k�����0�>��vK�L� 6
X�<	&�Ʒ���'S�(�	�m�s�$��N��6!���\��3���1��@��PN+'��������S)��������d��.�;Q��"�;�F$��C�4�X��3�����@�ݧ�!bG�0��\4T-�w�Dp��9Rxo0�e	H��ۓ���L�$O#��<��;���q'ع�!�=Vq`������`����t�'���J��.���@
���c��CX�lW��=^��v��zt� c��E���Rw��:�be5�YT�p�|W$,��?L��m�tIC;�"�'�ErXЁ�d�F�,��x��X����6M|�?L�\�]�[���o��G�v��g�#/����y(2�y��d#���?��{5�������:����g>t#к�G[�n�"R8���[!��%��E��of�3'�OC���]=+��BtXq����!R2���������|-�����\�E�@�jW�6�ɋ��1������9䷜��O���@�6���f�����~b:@]���)c��ۜX��S
"n)l��:����yyq�ढ{�U62Ӭ�[u��0�.�C�E��E;hO��S2�D�ڜ�������a�w��{V��D���vj@�ڊ��Ny"��c8� W���ɣ˦�k����"�{�����0f��Zw<��__��x)�v~�vƂk�4`9�N���#Ԝ ���<�� d}]3�����%��}�@[q�t+���Vw�JJ�����H�e�t���1g�ɪe����PU�:GTO���L"��l��47�N%��o步'����|�\ٯ��1�N��k�?e��R��6苂Y���z�n"����������8�#��S�^�,=D��$_�*��Ù�����I ��?�~��
;y���o��<\v�|	mђA�R��$��������v|���ôM���k;r� B4%�xhE�X1(�T��U��?��ڷ�%Ԡ���k���(�^��>�Z�� )ۗ��ڪ���v-��Rp?0=Ń�ފ.��r炆.�/'TH�x��>F,�n��z[��5��G����f�]BoLUW�")���C��)�]�?pv3����9���jA`����8�qtC2��_��Z%�T�^ﰅ(�6����fnm}ӈ,d�S�!с�㚴�����"$��-�WYb3V �	̲i������~�Obgn�5���LV�*A��Z��h���-�SFh���L$�y�>�}+�7�&IT��ޥ�
=��d�7a�aT�(�x�~'�����L����ĕ9�0j�V]ef<�i��'�:�4h`��i�m�Ǟ��ȩ�?��F0�K�Q�?5%��.����(�f���������l8�A�md3J@��H?����;�u+����������;�&{^�gM��B�"�Ǫ;f��yW0]�ʢm��]R�1M5��*RV�.���&1�r뺸�Vm�6�z簦|oa�9{�����^V]���]��7�/�M'�/+u����`���VBp:� k���mo�sE����q�ô%7�t����o$�'$�[b� *i�4�$�I |y��`�ˀ7p�R�'�v�H���ư�%v(6��ud��3�]j���Z�j�;ǘ���,:|��jv����Imo6�ߴ�j��{�W�.���8�$7Px��rB�h���]2长�u��Am���gUm�!n���7�Ƴ��vi�WTR�3�=8�0��ϰ��ˡe4}L��~mB�ޡ��hl��^A�ڸ����g�� �;�r](x���䨜$��m�����_F�7:��9P����GM.�R�|�c~0z!Nyp�@�ŕty�u ^��]K]�Ȧ�.c�O�D;��32D�7��[Pho
�K!3�؞���Ol)Xsm���o��XOX�qPZ�gx�{�M<�4d|�(&_�g����PFs�+��f?�Fd�.�-.��v�� �+ �{�W���پ���{�*Ck����#��A;_	�,��}F�퇻4/���U����01�M&�n�B���w�!ކ}f�oB�ư
�h��)1:m�*��O5a�1���hUZ�}=����s{����;�0-�G��[-x�PS"��3���U�g#�=kpղ�+,�,k��ϞI���'즇��w����X���-�c&a�l���%�7jW�=�x_�E�5q�E9F��w�&Q�Y<_k�D!��Q��D;�� ��|����U���L�@@��2:9�[�2�E�!!��%L�����]M'2)����A�ѫ�>\�R�k�E��,�|�zV���{�����X���Vql�SE_�LZk�o��S��z���q�bN,D_����сJK����A��tS2V}�섆a_7LjE��`�0r�Y��%6s�Gң� vUI9=A2�bC�HIߢ�پFa�Je��՜N�jAbN�����ڰi�E;Dl2�t��N�,����j:�$��;�k�8�e���<l����%�A��B>� ���$�Q�uk�3P3���y���z��C��z�h柩_8���+����$
���+������W(rR�IW�	���{���X��^ݜQ${���0 ������諏]�^�<�M���S�����:�zF$�l�[)�[�P�a�@��xh$5S�g�4��,4(�
kN'�l�  Ty=� `�4�f
���P���N%*v�z:wJ�E!%IUxK��@J���H��H�ے�_���A��dyt�Ѫ�*��7�f�9�1Q�E��tV}��58W���:R#�)@�F���S4E����qJmт�V�RVA�d�T0� ��?Tʗ�:T��a�^'���j�^1���Fl��]x}�t�	}�T���c\k��%��9�*qK<N�#s]���j��%�qSO���������g���05
�	W^��R�4K�-sik�M&�]r�l������j��=�b,37��.�4�}�_ym	1&�+�5ziH��,��?*�H+��m$5�" �x-��	����2�����%饽ƇUi�%.V�~9�/�g 蘴���1����.���7��vM��*@p��t��tE-��-� S������E�%%� 5�o��\�E��Q6�P�(>�U;�V�<��<�]g��8L����ڃiM1p6W�6��Fq��a^a@U�`�XՏD��{���D?�l|�P1��P�^6PkK
� #2�1=�w�j�k���w�T�D�Yו�+����s�������G�S� y%J3�c$�6�Εr&tJ��R!�ȡ��\ihH�	�Q�GB&�-��S�X1u�ۢ�����a��#��0�sP�S���99=K��(/xt�y,p�]+��:�_���)��;����\Ʉ��޻$\;�>�;�̘�6ӭ��j��Wϳ�:���'���'�yW}��P�6��@<,� 5[ل����Q��Qy������%@N\�=�e�rN"����_�Vq�\b��!(��.�A�zpO�*�4v�
8k�L�7����	͉����g��Ec��c���n�M��V��-W&��,��/~ɑ���OSp��HMp�)�uU��;m�7w3���G�)����+si�����k!�^Y�}̲��#h�L>�cYjFQ2���v��@W<O��I&��?,!���.�g� ��v��|j��ۘڿ��܊j�	ذD��u�8�u���Iɦ�ЮdT���Y��Օ�S�ϰ�~�6a����*�ZROJ�"Xc�'~ygR2'7�0�Ysy����Y��3��`ꩻ�Mл��Z���	9��@T�n$�NN��M4@-��w8��95I�?6��h�v�Θ�T��(����]��Oligy�=��
uR�fV�]*��Pi	�G�F�k%-Eky8>8)�.���P�+	D���F;x9��9��t��:��#:`�B��1!��K��˨��f�6O��/VZ:S!}m�[�9����e#��d�G}-���Z%���"ɇ�p��h���&.�B�t��N�|��m�-�S�����B'l��s��)���RI`�zӺ�Y�Ac�]&����p�}-���!�Kڟz�N�d�Xwd:�՚P�s$)�Usi�rJa��]��Q�e���j�`� o@�s�t��>Q�yO�6�����d�+}�%e�,jD~,v��9_m�8S���%5h��P��˾� |5���};:��M��腿T�9�G|�7R��-��t��?�ݢa�����w��1��Y�� �}|:��	�#�U�S\�Df��
w��>�<�9N���(�
�����l�h|�H�C��n���զ���P��6RV��Ͷ�A6�J�� ���Q WTu�C�~��;|�;.��Ԁ�7�y<������x�ʄnj��*�q��/����r�#M�1[k
��:�ϵ7D.Ws��t�YS���k�)�����ns8��=�'�/��i�8H�`Z�W�}�0!�.x�����d��9�I�
ŜO\n�.�EvV�he�S+�Űa@�}��F�f ������M�E��������u	(���&ڡ;UE�+��/�a�3��"���V6f8X��L�;ݛB��ʙ��CS�HaͲ�@#m>�(��A�t����Q��Nх.��9
�B�8��W���_�s��S��͍a��6�چ��P��-u<� n 2v\��--|bH���]YknQQ�V�X�d���:��F $PA�.S���؛G3�o��{,N�W�dh[i�M)�;�X�h�^eo�%�*1z`jf�R(�����B/��d��@R�ED��4���y�e��-Q(eI��Ml+>n���\r�;wzd+��qS{9�7�aF����f	�BEOS��*'<�G<�K����z���"evFi�1t��q��<������*��������`�Yq�@m�|���]e���R��s�Ȓ|�m�UE�����O�r����yW�
����)b)���hl,3����a�&�1�67G�Q��$	*��
S;�� ~h)��E�@k9P�z?1�VГj��ިy3�H�{�yGJ����x5ޘ����Ô���X�t��Q�O'�M[���	5@=zf�&cǺ���F[e���7�³9�4Q��Ͳ�le�H�C��#��M4�h�ˢy
�~�}h�r�z���7���G+��,�$�V�t��V���i�s��Y}�ڶi�s������ǿ&5��!}Ŀo�^��+J6x��#K��ލ�u�
 ?�n5��et��xŝb?��%�bNPN��y���^��Z�˅ik�p���dB&.[�9g`�e�%�Z�r���ϖ
��z���S�>g�B�֤7畺��Kv/�Р�>�e'^W&��D���
��c.���3�2 '0ѐ���J�\�45M%K��+s�(�F�r]!��wc0_�at�r�Q��Zs�fI�g���.��a����ME�F+b�u��N�SWA
QOH�fx0Fr(�yy�-\�V�2��)��0��2g�)�mJG�k(���̈́��t��^�b2f Z}�ߣ�|����F_������� ��y4�,z�^�ǟ'��ğv2ʁ���g�^E���;�A��U��ح�릗k{��S��?��|]@N����x�U�Ɨ0�YT ����7cf��%���yU�a�l�C
��������˽�_�v�֟pp��	!��bM7�\w\N���j})��r~����أ�}c#+��G��o���f�d<���e3�+�7T��$2}��>��k�����^��V�G>����	f6+�����Ź0 <䅇��xgؕc]][�kE�a��v�V�|^LZh��=�-E+/���!&R)�\"2r�L�d)�m�䭿��������v ��J�P)WKkF���wim�R���fȱl�V�T�R<�V[� >��K� �xC��淶� �:)�>�x� ��Y�,�[w\{�=R�����&������:<�;��Jo���#�`����4����x+<����J�x5�WP9�l��O'n��۪OΓ�LP�pi�Æ;^��p�7�`:[��̣����58Oh�����KO�%�&EZD�а���ū��N�W7�[%fW��]v[6�Jp,? ����y��)�.;:Om�;?Y�2����p���l@�ӕ�M������0�}�A\��&}�Wjm�߬�t�w�[�/����+� �ՐiuhE������|�A{���Z8�Ng���jеZQ�H
�m�y���ζ��{�@7+0$�1��}t b|4Ȝ�ػ�Ƥ�p���Z��L5/yɄ���_�@�z�����	�;L�w��W�Ez2�2����F�Z��L-IS�T��4n8��	�Z�3 ��ތ"�n���,�)�]������	JS��Y�*7n�۾�+13�_TX?s��$vu�:�����g��a����:�T�57p�?�� `�.��Ը�ݴ�z�f8څ�>Г��P�)t��q,�!�[5|_J9���Y��u�N��D��'�x�D(G��7c�n�5b,��|�+a��?��
�
�.>��.a����d��B編y*n�z���.
QLpMkHZ'�2�G'���Q@�FcB4�:��������9-u�qFTHq�S�+G13���6n���$�֋��W4�<��J/���y��XV�h"���7��J������n�ܚ����U����[��}ʘi���k�Nny�͟��d���{�ӀoM��Z�Ŗ#�}��A�0��5� h���W����D�V�Jl��襚mR?�0=�9v����]���U�"���#n~����7`W� u ��� �T3�	���_�Y��D\�&2�8!֏{��1�h��8��g�ZRd�ո��c�A3A�bt�v����u�[X	\���PIM��˧����z�t��C�_AYuB�+?�m��ؠE�R0MQ7�X������C��ڈ��&��Q��4�E�g1�t@e �t.�%G�@G��Fa#��#款�| �-6E#c /^B�cb�?j��2)���j�D�^�J��/CQ�ƻ��68E�?�>�N�$C���8��'�Ck��x�6��:����"��<�u����J}h5�c������T� �2�i/����=T7(
�:� ��%�y����Z�֊$���.�"��G4b����v� U,�3�J&J��I#s}Rh��:��E_��ֵ��0��J敓�A�Âɘ��_���ް*�L�~�FPtf�"F���.�K�-�d���U�����7��Ha3�z��X)5|=
\���
�� �6R�J/�9B�*�O��ي��V9Ө&�#:����\�n�@�"��N<tR�J>����H.�6���y�d¯�]��V�����o.���4s I%o��زB�}�8
ԐiK�.l���N���h6�3����]�e�oRD��@���wً%l�:&uR��p]��Xl��A��*�F������8�y��('b,C�<F�I�pȜ'�L ����0ig�~_,����=i�^�wr{����VΦ #������tD����M濮�U/�"-��9�O���P����f��M�x�v�7z���Yפv�RT�^��m��5,��h$7�5�p�{"X�`&~��)��t,�O}t��ɀ�a�퐋3ٍF[���g�vE]��B�q\﯀�	;Ńb��|w4�\������w�+�l�_��ж��̨�1d>M��p���0bh�0o�H��j��O�2�d�.�����9��W��!Y��v�%|4Y|�˛�s 4T[4uO dΓO�'�'@[,Dp���zs����L�x���ԩ��"'O.@[��J��m��^���vӭ���������p5y����Ė?���Z3Kc#NJ�ͩ}��f)ы�+��2އ�U��#6��*�7Ĕ_�|�柊 ]c�\el��� ��{Z��rrFh3)(�����s6�����R��<#~��X�c`��Lb�C�a\P�����*'x�Ӹ����gu�Y:�e�/֌���hk�}��׭���4sӂ]ʿ�z��nE��H_lE�v{X�a�P,���RJzI͟�OD�f���*�T�9��ї�i bF5A��RL��d�A����ɇ�W%^ll�r$B��N�������é*�Jf��!e�qΗ�,�0R�(
2��(1
�nc�Y���{ɁĞ��7�	z�}}�/y)'�\����9�a��t̑�=
�"jx���M���r9���[�w!x�} ���U�v�.�E�%T�1\e�?.�ig��X�
/�и�����o�\�hoVA����_sGT����n���w迬Q�&On�9ڲo�ͪ���u�6�"����Y�tH�0o��G�ؗ8C��mxi^ۡ�̮GG�����	Fi#NY����(�bw<�@T�<�N�$0�c��?Z=�y�M��+8�+��+R9�
פ���,q�O���H��wʭ����8� J�@�~���z��7�oA��˘�ȅ�yN�͝�f���;wcL&^�C�DNs����,�&���~�ޓՋ'"z��i�0�U4�L��J���|4rM@굿|8^^�-���Γ��_���/���pg�l��[ �4^yC=@�xcj���l�5Ԙ�����O�O�џ�E���Ӟ�4�%�=:�8����4��-�D�$H˒dhCo=�S���,�!���?�aB�T�F�	����`���nb��,��:��ü��<Ԛx����c�p?=HO(�"|Ƭ��z�ߣ���\�]��Z9����u�4Rf:˱Y�� ��A]*�������
2�-9q�Wu��o�]���&�W�����Gc�Β�d���H��s�VRwI���=dNA�TѢ\s����	 �<q��U��1�ΰ��\��`���N��A�����N-�eߜ��u&˼޼�0Fd����������+9^}���
��5f��)�����E���T���{>��x *K��6�|!]�'�j�_E�nk��`����k�9o�0���P��nWS���_%�WR �K{&@�L6��:��G��('7�m�eT�U�M��`�sU����e���|�#��7`��]�V�M�{e�����HC�0�շ�X(saԖ6}����i5"k�|y�A�-�2��.���2\�[���ْ�#�$M�ϛ�)5��Te�0�������䖼�HM�⇲s�a*��nv8�<,�D�*
F�Hu@|�"2�^)�[wq.F�ey�Y�-"A�.jr�h��rw��<�����w��ZC�❩��0V*��׏�O��z�F�
�J{���6"������L��2�zX�y�4���7[�����j��܃Kw��n�,��,�Z���f�d5J�����!�Pz_��s"'�bgH΅ҵX��qp��ʹ����b29��OM���%ր�A٨�N���Ԅld/ҩ�D�U1g��eO�8Bh ����Ԝ[ �C�/�uuN3.��Ӗ3���L�do��U>�ˬZ�r��*����P��j��.��x���"�� i��ai+D��>ph�̜n����rX� _~�z]x�X�?�)����� �M1���t�$��.����k� ]>�A�#l;��:n���t-'�ý��ˆ3�ɻ�b�&��i޹�.Z ԍ�$�>�ئ|;�Uh�X1]n�C�y����kY���e��K��Z��c����⎄��S�8��}�9���r����v��w�����]K��IF��- 3|iz�O�6I	�b�xx�#"��P���#�w���+�FXb)�±W$/�]i#`zW�5)�o���^�u��18SIdYW�r�A������c:���y�ќY����W$��I�.������B5����^ώ9[ʜ���w'��w���g������~gT؀��8��yS���JX �P�FYl&!j�W�ص.�1�E�|��*i�Uv��y^M� [�������t��+$f�h�d��
��V�ј�H��բ7z!�vF/����( 녉<�MD��#�C�_@�mP�p�\a�J܆��l�.�1&J�>Y�F�J�s��w a+*;,gh��f��Bb�j���#�T	P6Jdo.F{jq&V�
�����"��2��"or�n�U: j�#�r�
��6�KLVM�aW��z���{��3�{��*h3*��G�ެڏT�R�����켏�*.uZ;S�=qb��02t-	�++��I�ݪN��_(_�(pɕ��=#N�JD���0��@�O�)�cW��[�=�J��`׃��^x� ��ҫ^�[~�L(�埌ܭ�����:��8�*L�'����C��C�Z�}"--!0�����	<{J�F��2Q9P�ղ�D�9����DWu��p!cZ���C*��%�ו�G=L_9a�+d(߭g�:S�)����U���=�nC�t��'����M�_Oc����{�������uZ�*a-�Ҵ���v�y��ho�/N���֡mC�3�E�_,���.��)n��gD/������M����ܳ��GCp��"�o�����V��P\��Q(;�����Z�O(�=���'��6+.�3���uW~���P��t�<��Vx7�2���Q��N �����s��ǙJ')H�����:`
����"5�+���Q����@�~�Z���[t�:���2a���b�\����6:-�� ��ɒ��:(�� X~!�(
�O.��������n�љ�4�����nAP�x��O�3�7���ag&��1/� �߬�LC:��C�����_�X�2�+�sʚ2U/I������v瑢�Jr�FZ4���m۠���:&���d��o������a��_�4��`��(."b�v�8p�����aE�<���\�$ ��>v�T�Zf�A/���#	�y��	a����]�l�%��&3���S�$�4R����D;��?Q�L���ۤ��UV�C��i�����l���!���i:�Bx��9�|��.�0c+|�@�+�o���.�(�6( �c�8�P�hR�n'�*05�ߘ�:�p��h��������9xs55Dj����F��ɰt鮆��'��οN�Kӓ�7�V�*>�|�ܞ�~��Ol5����*�y���>l#h���^H�\`�p���0k-.h�Z���zTy�)�0R��˽ ����/�+�w��ϑos5&�Ψ�����$(� �28P�Nt��q�N�ڒU�K�&]a�(X�P�u�HZG43ئ�C]O�Mݏ���UƩ��V�	0��	��<Cdd�%Ɋc����H�/{��*�n9�1:j��	긍�}�VH*���Q�,p��tP���z
L� �֑�*^�(��g0gu(;v8�0&c�b#����������HK��'�)�h״,����4}uP���>R��R�%-����~3�O'h��p �R�p@�\���\�'hC�����[�����:P����g�I�7t=���q�^��DU��o=�Ow+�%p�TV��O��i/����6�*V��b�ϣ
XP8�K��n��}K,"�2����i�rJ�2��S⪮�c�'�ŷ�y�G�I�����z�z�J����}���v@P���-ko�ÜZ����ap�l��ًo���sXl4eUZb�����g.�����]�/}�YZ_�_$�H�<QH���K?�!�U���
#��9CA������06���}8�Lqؐ]����P,Z=y��,�� �x�M��3u`02�n�6|pgE��	��]��Hv��z�_N��B׵i�R�l��ӤOP	`f$�vA/�Z��e<�k�J���"=ȴ�*�ʌ�Q��'��x���(�%^�<}��_S}�P,V!~�t.�2���Ơ~f�X���ɘ��jN){�p!�MT�����%=����E��C��#�y~��-�dt	�*r)/k]�#	|e
铏�:��4]R�$����~�z�kF�X'�a�����"e&>h�����_Y��^�j���L�,@�[��<�4� ]��t��vF�|��=�U]����C��΃���ٜ
��`]ܬ?x�Dh�*{)�7��H$��v�����X�#��fb��5���62-�ѩ� &��٭��4��H�j�d�2���<��HY6�
"ȿ�����5��K��JD�%�?��N�C������]7^S�j�_1&�b��z�wܽ]��7�F��6
�i�21���EW�o��/Q�I�@HF��,��1g��DV�e�j��<.c�?g���{s¶[�-����es�!q�ҰF��T�g2����f���~�r�T�Ԗp�eI�]!y��ICDh�zA}�g���O�5	P�V����db��%8������<c8�r#�J��{S_s�\����;���J%(��5���h,5]2	���Q@��V��2C�V��@5M2/2̨5��}���[����ڡL:"��%��P�Z��������R�e����f�E���56G|�Y�]�m�Z�z�/��nM=��A�B�T�������y_mRi����(��+)$�߰~��� �F ��h���j���ρ������_���D��4��
�G��ސ=[r�#���L��p��/��<ǿ�)�i[F�č�o�?�����/j�͠/��DK=k����������ñۺS�Z��NF�
0*�0�J籝��I�Ckʗ��+�V����)s��`�@��4��m!'���S�'�	Ҏ�{�WI'��e��c�D���a�i���X}:��u�R����|�ڎ��<G�|�GS&��reW�AaN�������Ci�^��t��fޢ�g����T��3�tCK@���]�����H㽜&4��hN�'Me K���?�A��W3��q���C��'��'�>�XF�n����o  �G�ng�n!H3r�F��p��f��������MP]��� "�	��u<F�5;Z���r$�|��ɲt�>��N!���g���o�i�qvϮ���LȔ�V��
���+`�A��I%+G� )�Ri�i;W�Tx����f�FKD���zM�<pJ�)�S2'`XX�mo�-ĭ�.�Y���82�YvL��&�g��.N����L�W�r�T���w�;4�%�;I�D�.�b��hy_����|6���7��l�u�Yj���S�Ν��r�6��G>T�Un}!bW�¸IUЌe�"}�TP�&�7J�@�"T�;7�S�)u�'H+�[U�Шp�#�ihTd�˄�[��e9Z6�T?��i,�ԇ��,����A��z�a�q���BWS����v
78w�U�V�}v�B�r�*��܈����52���������Rr�w����rf��Q}?�э׻	֖ϗ{��,"0K%��];�n�.s�EWM�5����0D��pT>�o!1�1;(�B;�"�W�,�(㭬��n0P�:+#�@�FB������#�
%%���B���ף�q�*�+��N���Ky�{}�+��"׫�/_bHPb��|vw�������X+�Sjiw�@H"��>�V����훉�FX7�)����E
TU�r')A��F���q�f5�x8kB��g�;��4��GXPIe�T��8��I��!�Iy��Z������y{⺍}g/c7{@�VlK>���Ģ�^lvD�G@���S��ę�ԃx�P���X�e� $N��+��¾7d�/�AV��_���4G=U��BM;Ř]{s�?h4�?k;G��7�6��#C͏>}!�����#QI�8�摣�,�
I}�Qȃ��pi��˴�V�!��!T\�I�G�s�����u�dg�3�H�ݖc7�X��ˠ����R���z(^%�,����YsP�w��/Bn{�z{�qm�ϔ�]R�'����@�������EF6U�B��@:�3�zd'`glKD�@;&�r�׷��뺚�W�z����\�v6HbTP�3�5����Db��	�^���Q~|'i(��Ϥ�N!�m�O;����J���l�#�.�1�����+�#��;v#�b��g����P�q$f��]��hP��]��,�1[��-S�\�H�
��b�]��d���@������+`�DO�)���dIgV����}�����}��jQD�����Ǽ�]m�Uu�/�3I&7��x�Z�<��g#x)���J����
��+�ԍ�gA@ԟf�|�,�S��ɫP^ֺ�x�8[��Ztd��%0|��ڀBGL	�nG�%������n�a8�tӔ�֣��G)��f�5��݋�F�+�?�����`c��q&ׄ�"��/��v�$�X=W��!��I%&h�I\F�Օ�a��fs�M�:I�>9�G��] ]Zs�Ǭ*�#�����yw�G&6�6�?�nV�1V��T{?���jͱ2�h73[�ҵ�@qS����Ų��&�M�8�QC�쓛�I �@\���KyÇF���p��i6���6
�e�.�o�M�
�i'k�K}��g�HM����V].��W��_���fH3��ےm_�~�~JJ�C��-��ߌRkӂ��e���G��1VD]�ô��nw���1e�܊v9SS��M`��8و}���T��V#�-�	?�$��+�؅�����_��J������v�	G?(n�q�	q�4�e�&��)�(���r\��Y8:~���2hJG��+7ۀZ��]�
��8F��8���c��d��T�HI��TxnB��O@����%�t����:]�`�[�0j)��_���MZ��$����1-����6��U9켑�,��P��6�?��-}��rMx�#�V���9C,����6zx.)����v��B��s���*2�^���N� 	a�1@�~���ײ�:@�b�?���� �vF,4��t.����P���H��5�b߭�]7A*r��O9���>m?��S՝� ��j�|%Af�c�!�U2W�r�|����nr?C��Q�ZA��a\7��5�����M�Oю�B=Jl����n,㴊�
T�v�=���W�-����|_�ly}S-���Zj�,nM� ��܄��i�&<�h�n�`�4�)�[�f.6���u2� �;-�9�;a'�Hk�rn�^�A��̵�G��ȱ��9lP�98��p�{P!c���H�}C~bMl�S�N)��2����/��?%	�#�yS��|<��|�~�$g���U����b�8c�~��=�(���K���l��Z>����	�Ƹ�]5�|���Nx!gAPa¨p���j6�J'hI&��c2�ͩw�����[Y�D�:��{�Et�	0����q	���h@�bu?߲����*2�9���������,g��[uﾜ�>�Xw�A�U��������L(��a�i�]E�XcD@��9��&�����NEg�G��N��W��TqL����9�Q>�ZI����P�KvMz*���pć)�d�쾊��v�b^�d=u��L�'7BD��Ey1�� �?G��1�X:��Y��f�B�ڪcDl�/)�������gYW-�=��9t�	�� ܩ�9:_���X�IĜ�����K��W�b� :�"��'����:E~���F�֬8����AL�8���U՝J/�*�<�_-��9L�X:�`����+#�S W���7Yi�B�5�od����mL�#�;����%�;L���Ѻ؁e�-��>I>��m=F���[j������V�d�#������*^J�נ��́�Q�� ����`���6�6��H:H���e۸�ܻ�E�щ��@j�5�ث�]�J�=��c��T �����)]�� ,���@߷��ӫ���:Η{���)��!k���p���[x$W Q�~�n�����-x�Z����L�3	TO�V�k|�2�_:�ʪȻ�y$�&o�1{�6�
�*��F1T#f���o��1����@������s�N��e�S9۞�`"˯o(��#��Q��o��bTt�,̧��jMil���`9��O�I����$UV���x�$M�D��	MQOi��(����v��m�@"�ʫz�h�^��gY��qԐ9���\�<�Ҽ�߲d�ڹa��6,sDt�	z��#s;��\��Dr�e��v�e��u-�l��(|]�&?����P�"�����(yԒǛ-Y��^)�]��=z���"3h��L�!���9"���@5����1u������+�c��dGA Y`�8�sa����'Z]n���7Q��i%N#)���f��G���F�Z�Yݪ�\x"O����AոR�y%����E�
Ø�OK�-�^ZqYXS���h\%�ߔ�)��q
{z��-len���'�����l\��s��"L���T,�C�.G�-�j�{�VZ�N(�ߤM� �x�֥��-����<4Y���ƕt��/���L�|��a��	YO(:;��rd��ĥ���S�����P��8a�x�������C�1�Z;ti1�J�	�9Jo�%fH���lne�Wa䧨�d�C���g6ʋ��;�]`��>&��պ�`�I������1��&�}��o�%�-C�_���&�E)N?C|�m��d���Az�^=�E	=F��w�Ub}ܾťV7N���r��bc�}"kH����wU'[�L�Y�F�#e��Z �3�4��n;�R�Xh�]��F��T�t�)��v*kg8������L���@/U=~�,sS�M��E�PuK�N�4u�%E���)��0RD'�2�r� w�ynGq��� kS�=\_�b�J�A��q��l�F���Ҥ��@=A�5	�~9����ds
�C2� R�Y��[���^~�K��	qD�rw�G[0����:I��f��r�m�4�uG1s�3�G�i�Pöǟq�g��D�o�
����x�d��l�d��EZ~i~<?��*b!�ZNE��3���.`��%����|<e����_|���h:O���t�����
�b��'6I�+�I)
�Z"�:�w�@�E��o���ܔ낻GΝC�_W�u߸��cϝ8���5ҠV׸�s�B�Y~�h�G�F��Ⱥ� �~�0cU��������E�+gc�&4�QJ�ȹG�H���=Q'���&�o�)��f�JV�rw��kjׅw{�{b+0��80ڰ������7U�2:����e�?����p�^4F��ȒՇO�,����M)��+NN�������b�gj�8��̋,+Igy2���3��~U@�rUֿ )?�>{R�T+iP�O'5�_�N�ģul�a����pLz���({�?Τ{���V��Voc�C� �Z���i�F^&i��HH݌�.���F/�|T�^�_��2X���?�Rứ.sPg�s�{�k�w~`���}�T����d�+��е2�� i/$�ߕ|	��E�U�9�<� ��x I��M����z��P��$iJ^�:݈�԰�� d�r<��#B�� �=���D��\\bO�����5�P�ī">��m]���5y�X@D����r3�Zv��Wif^��A$	��������0]Gc���ǙM�����l�ߪǯ�E~��8a?��<��ZT;� ����߮M��8||�o에4��7��t�/�*�$n��cu��]�����
$�E΋��{��-ҲD9�RJ��fqW��Ӥ�ip|��ݕw��x�Hͩ�WQ��&�^�?�b��$���lb�ca�Jƃ�Yп(°���%6�����~<C��#f�K��[�|(pa��I�YAҗ�Gi�ö�� 
b�Bp����~�,,'���\"���
���6|�(,��a�1an��7D����)���ܫ��T��O9KP�n���:��� f���WE�5o�J�QB��|���]r�{ ��dO'���<�c��f=��e�`d�t+^��C ���p�9��4���y�l*��\�LKgU��id���ʅNׇ$��pf�[�-{��l˂yJ/�*E�!�e����b�����٫�H��H4�yG��g��I�+��{zy�_+�)"�;��3/�hQH���ީ���t�:Yu���u���*5s`��D�f�v��E�%�͍K���=��[n����ˁ������ֽ�)��A�Ζn	O��4o��bf��
_�v���*<�X��[��n4��(w�8�fĎODw_���O�H���?��nb�n�f�n��^��ǭC�ޖ~�ny�nrE`���x
�A�ܝS
ޯd��f&�������u��w�Z����~�z_���gi[�N���0�9Ì�_�|�Tg�xn��UJ�`�C:"��WSN	��a�S���VHw~ ��T�����V�G��_��%�xT�m�j�=Y�}��ۡ7�񧗤����6I#�o��������G��� �AX6��b��(֠�ϲ���toUQ�@?�rZ� �5�#D�M���H�4�OW}8ܫ��n�����(d;��͡S~l �z����ۂ�x��i�bd�;(B���h�.�F�
�_	r��l��1L��.��+�.�B��!Iu/�̙3���me��ȡZ����?��Ӌڐ�G�NR�`�{~�$���!�ݏ�{�@~&�1j�O@��r���FIŮ{_�c��	�T�?�j�H������3��_/�K"�i��1SC�u�q���E������=k^��W4t�kW�`�|�}�Ǳ�����0EMvޡ���g��%�ٝ���L�T�#qYoQ)�e��)7;�lXx`"I��#_�N�p����dH��!T���~�A�J�`�������Q�k^>��<�()j�6��Յ������>+�et�.�x�T-nqdݣq����;A&�wm���@MJ�ߞ5,��a�മ+)7��BJS�;�΢��$wp>xS��j�)����t�/}֍u�0j���/��
1��F����F�M��G!�v}�;U�����8��H�9��L�@�҄V�g'n}��I�=��w٥q��i�'t�|`�y`4��꘿������.cq��y���	��et����-c���Q9Yp�������|W��2xzRp�C�^����y�RA�;~�,�Ww�-�ZudY��y*{����[����&AR����F�����H���>�	1ZY���j����r|�c��{�6�#�|��٧m�i.nt���X��|�����כ��(���n���:� ˇ��y�����_�X�o?y�c$��L�P��Kx�i'*:��$��63�#�R�����Vp�!��ȏME���w�`�t��$f���� ?�+�4òE�����������>��)�H�0^�������\�q��ȭ�e �����ų�g
x׎�8=S= ���ō��]���:����=��!f�W��;dOu�	�1��������BT� �t		'�̭b�J�U�+����?���94�D@R�4v�f��r1j��q�`�٣",�P>��ee2����Ļ�,�ܹ��>�Ù�~�vc:�xSF��E���Y���]jݷ�J��9�;;E������Q�CW�k�S��w���;�-�����>3��J�J�.����{���}y�B�n�;��t�:���g��VW���wk|1���Y�2�iF7�wdY�E���s�R�}aN�9#�m����s=�Hb!Ɗ;[�ckr`ǌ��'��T�S���#�!�$�B�x�05>2bk���4�a���<�6��4�2-pS�W���@���wN��YIP�\#h����e� �c���-�5�?����\���l�Y^�����V;�d�gE� �%'L�r�d�^f�U��vrF�	,$�I�XC�6�l4���t8����H��X��v�n��u8U7�Ǹ��=J��5���
.�r-�j��1��P�sr��g.M-\CRy����2e��s2��\���:���l�cf��k���
�z|�4K�\�� ���'Z6�S�ƳC���̘*u8�4�3����\��ZX�cF^����H^�x��G�y ^��hTq��A���%����q���/<' T�j)����QnW�5�DՅ�$���&w�U�M�TE�-�[�$�i�."rTmh�r�M���c2���w�Q�"�Lő�w�\8�fn�!���a��]_[p�
C�<��u�t�r���+�,pqP�M�% �_0�� ���G>�I":�:g���4њ�NB>eGN���v`��TD�rN]�����~�oK�3��C�uȁV�f
�̼o7��`Ʀt�a�^E�v4A�XX{�6���`��h5�h�A��z�;�>�?F�2����;���_��y�#����
J{�tJ^�a��7t���H��c�H��J��-q`��&x3ŊI�5>��̻d�?���r��ǘ�^v��m/��cDA��m�"6P��餴����%��@p��
Ld�g��4���#:-5��>!|�I\`v�e��hY�`N��22��3�ǅ�R�B{Ͻ�4��%��,�yTפ��]oxq�����p>!��BI�ȟ<�)��?3�KD��|���c��L�V'ey�/�T-^�}��fnH퟼To����䟼�" ��W����7�p�E���ڪ���~���_�kp�@EEݬ����I=������M;��T-�E�`0�p�yCױ+O��Oܨ�@�r��ǒT�WbTCR-3}��PhZb5��h��Q�0o�������b]�(� ���z���Y�dȜ:r�)��Ӯ�*-`���l�Ti
C53xh�F�YOC<	���0G�hq���I�68
P�l�ˏ�+��>��ʇʼU��jAr-V��L6(�IrZLGs�:�k�_����f�V��\*e+@�?�=��Ĉ�H� �;���U�.��xve�L�[�H�Qك�~�S���?��6�/k/n��wȫ�><ܸ�E�������/��%�'��j�h6���t��<�o��+m����la��|��Ѡ[�L���qLM���C�I]j74f����P�,ﮭɧr&8e1o Ϳ2�L�!�=�����Ԕ�E.צ��%�gjmR4���e��#�Z-ȼ<�3�f�f;�����)G@9�����Cy����g-��<N�f�������*�O��L/����oQc��KU ��g�6���[����I$�����ݫG��".�I���ь�l�U�7��\Ҋp��|�>Q)~
���n
�>���37e��ý"*�I����}g��p�j콮�>�Z�(~��'��ȤO�`K�)�ޔϑ�I��#�� �.#R�����r�"�jq���fي��������q��#��.�T��R�r�?�O3��c 'D����o�b������E�(� ��RM��Is���9X����O��[
,������~����l�x�+��\��e�εkK����	�ʿ�5��Vu��%���Ϫ>u2��
Fڹ�r���y�RA_U*H�$+r�Z�n��*��a�]�(�}�}p�Q~Vԉ�IK>B�����f� �Qi��oB�����5���,knD�Yg�Tb��HŲU�GD�I�_�"�>�-8ؽ��ͥ��|LFLD?&���쪣$T�s�,ۋUU����T"�"�Z[#0�1Ә�6Cҷf-����Q9�QeV���9��z�z$�#	�i)|!S���!'2���1�_�K�FNW+J��� �-�#(������fN6 �*�nmP�������A���?��^�ԉ��f1w'��:)��D���sS\�@��M
�T�θfץ�bE�Ŋ���PGs�5��T���6
�Fn���_��64����~�����	f�u��D�h[��D�U?�����"S6ŀ��E���j��:�46���%�Jư?��;�����\��~�4�ɖ����TYw!T 4�u%��L�: u|��V�Ti!���Vx��cJR�F叁V���-�d3��8xl]ت��������f X��EYx(>��}��,}�1�'��/����=�PN�)��ڭ6V)��F�Yby����R���H|[���s��R)����ONe��<a������B�Ɍ��.%a��1���������zVM.�k��	#�r?QeM�w��"wզ����ϵ�FC��׎pu��Ȟ#;i�r07����@��b��SY���G`�[�j��Lp�%��˃Lv�XfS�R?���x�N�/L`����4t�Tbt������>���0@�����z��ij@��yrX����s�<ѥU�5��EC���p���	��{�+=�fڿ�W���o���	R�v9e�����VUk�.z��x��+^+
.�9]1^�b\��[,�g���5��$�	*�)��G�FJ��~�Ԉ��$�K� ��.��������}��_�w,�1"���k�14 Z��J�1�o�W��;l�܅Tŏm�"ǽ������ӇS?-O���kjr�H����_&��'Mn����䔘�@y��'�-7Gܣ���i��8	�����U-w�ǳ�4�	��$Ł'�(d �a�>�`L�5��4hq���mWrDp����1iR�8�M����vc�_�j�S��5+8���+	k.BA�5&"Y1��CM��~�����Go�~��J�L���P��$�T�1�WEJ��x��C20�;�5V�]��A�ט�����LpY��WR.c�'��̋!��/�1�3�*��/�	�w��lu��j/�UT>���Ȍ^�~/f����~RS�������
"W�6 ���{����U�s-�G����	8�D����	R�V��
�r���?f�%�rJ*��1�.�Tx��ZX��d��6���������S��`h��i�^T�Q)���C��i���pל��&�oY����%s,�4᳂�^��H��6�U�Y{�6!]ښ8�����)VW�P&�)��G/I*�NO�L�:�;-�DТ��UpZ���� ����%��?_�u��	#k��+�ߗ#������w].�s�E$pV�)R�~�Q������0�:ޱ[���\��V�;/��B��
D�G�7��_4x9#?<�%-!��0���@�mm�p�ԕ$'ֽ�K��	�4�:�.�VD|��/��<!H��Y%h ��=����2>�}kD��O��dz}�Ir��a����If��d� W�O�h>�l�f {��f=�݀�hX/���soq��1u�c;�i�V��j-�����6䬣q�d��#�c�~\�4oʉ�m���+��q��z0��b��F��]L��ȱp�~�����n~�8�W!�5�����K�M��j)>u7�IN��4ouE^J�'�Ճ�[��\m��G��]���!��h�Rg9�B�
��!Sr󚣧W�lX@���*�i�m�s�xNxY�����[�hQ�q��:�bh8yǜ<#'��}�_�Uߞ[��>/��ϴ$jIƺޭ��(Z�n�$�c��I�O��PiT�p���_F&i����c/�Y�>x�:*��'�ZV$0�2�ާuf.Cϟm�Pe3=?(?mҦ7�o쌲#�(�y�CΩ��D:��+�N��3a�!*N�l6�=. D5ih�j����-�uNJ.�wOg��R}�`]"N���O���\���P��k�~����}��
E�,l�n�~��(��ж�f��*���v�tys�}�N���ܤ^2Σ�.
�ʞ���N0��H��+�av�V�k�V��áw�����>�0a𿜤�] ��D?�oV��1�q�~�A��8���]��(�D���۳׌����{�Q�F�]�%��%4�׼�B)�����)#�_�YXºx���)�,~�j�5s��I��{u_�F �B\������`jetv�v��G|���Ԁ�Z�[g�7:��*�&G��XJ�l뎰�=�t��{)"of^�c$j���;s�{KN�䢾Ml��9rl�$�i�Bf��:c�L%^X�T�i��iT߳��_:�qq��~)Y!{�^_��8��Y���WLW[�e�-�D�Od�����eO�2���]2d���$ђ��+�X���խ�!���l�.���14�G�G���O���5R^H�\hp���)W\K�W0�1ÞJ���i��Q,x�߲}�D�s��zu� �9H�`т��=�8�0;'ݽ��v��3�b�� "(Ǜ��B��А�S���ܑ復�"�\�ƈ���>�d����[���k�<w$Tj9MGƹb�e���Ii�AK��mC�&����I�7�.�
�3�ጿ��:���~�?F�M*���9�hǧ������m�A7+��ɹ׀�V��ö�{*����1)�'Q��T��&a�b�����B����Y����@� q����]C�QT�ʫ��C� �����X�ٰ�f5���dU��p���E���c���&�� ��e���[S�6����g}����.���G�(���αY���|9c������*���zQDI|��ڟ���D�
X�����Qs%�9	�\�x"��O���U�>����fLT����±pe-�p��Yd`P�Ac������щ1}-��$W�L�SC��܏:?�`���e�/�V�j�5}u�y�3J=�~�HPG]�p$�wQ��f��to���\�ҕ��@W[��1�_4���X'E�a>�"�̹B��3���hI���,�2��l��$��y��Lj���&���P���B��0ҏ�35���I;O�9�S��Q���m�fUi�ˢ{���+���P�� �%�5�v!A��^ÅO�T�k��sq���FDZ輵�%���%�T�/x�Ob������N/e�t����U�5'Z�*�GɃ94��o�����d ��Z�/�ƶ�}�G�7c���:j������3�Ƅ���gh��O���j�&1c%^���p���l�BM�)���b�8Z4N���??0v�׻+C5K���������#���fB�8K�@B�(؟
�XC�)�ك:e�
����i�E���h�mH)���I��$���\<�WF�?�{�Ʋ�
iG�w�엪j��+2RA�S���UhT�X�����c͘����7r�h�{QP�EO���L@> (Vm������_���Ciz���u�5��r_���h������ȧpQs��g7��M�(>��ɷ��̺��)�?3����.���u<:!19֜��F�EOߓ��1k�H�g~-���
u�-����Y�ʱT���.��=R�F��{��1����U���q�2��_za�IIZ�j�p�"���I�n�ڷ��=Қ����˄)�g�4���߿6y%�7\(����|�D�Q�'V�%*P�a����`v]�:��N����Nʑ�bB�A������z��'ؐYE��Gx	\R�	�O���=��sd�|`��-��|�8�9R�}T.�Y�N����d3�A��X�c�Dm5(���Ǒ+��Y\o'��"��b�o�3Ps�"�d���.]�""I/�_���DR�i^@��1,ͬw;x�c�)�rI�Q�}�Q�C�m���g�:����:��#�Y1�k
HR���ߠ-P9B�nz��LUw="1?>*��6O���]waE�A���R��;�V�x6��Ge〒=�^:�s��.~k/_R�.�׸���E<
��'���[�N���7��uc�*J4iyº�&��՟:3����/�	&{�����	��}�4w�Ӱ�H<�m)��)��I�13����q�lu�}�.�沴�c�4j�����m�ov�l�{"�����4���0jɎ���kФ��B�m[�5���IRy6�^�Sv���9S�j`���:�.,�8��-W�*Ǒe�����IH�8��R�WF<ٝd���(���Px���]�:k+!��=�r;�k�#D�"�VKB���,�Q��������	J7�
���2.H�Ks�d���]X�j$Ak��*���W�OB7���[��p}A����PLy&�yv�l��ک1���	�G�wÅpT������%���-3A�BJ� �>��ij����j=<X H*l�A����@��jI{�V_�Ϻ���Z0��s3�����_�5"�G��җF��!����Ol�|Aj��[���w�O��0����"����K�P�mmiB�y7l��LH ��3�>T�\3v��w`�x�ß��������N�t�w�O�������at�����?6��kP=5ˠ��bUX.��$d��i�Gv�niI#�ꜻ���Oم�M8
%R�y' �·�����{�O�X՟��}��I2��g_�ȶ_�����ΠbF���b�j��v��\%�E�m��a���;V�[�j�B(�MbrO�.�̙cV�0���(0��B,�D�/]w��p��3/��8�v��E��3�B�]�r��^���<��U?r�V�WR�}
�l%��w�\P1Leg�s�eg�kg3��5���	�N��2؅��|a%�B�^p��	��ꃎ
�H��0�v���l�7��a�FˍW��6ʘ��k����%P�Vɟߨ��l�'��r�JʎS:8<�k!wl-�?�	��3 g��`�DX��ۍz�ah �C������B������|{Vfw혆;���2�2���k!��F=6���^YK�:��k�!w�g���O��6�x����#h�ܠ;㍈Ȑ��v�^��x��s!o�jv��l�p�2�2��ai�'�JK�h>)�(S09�����}�鏹`���]d�#������C��˰�N\��Al7��0a�����s-�r�b�x��ш���/�M8�
�RP�$j^	/�4$>X���@+��s�Q_Z� �}�7������N_��d"��7	w�|]x,(�[��4*kC�������B�����ʊ�d?�L�21U���ea���R|q�|�������+bi�9!��l���&��E�:58���v��Ƕ�ջ�L���H���0��kLb�F������l��K��0����4��ɭ���o��y}����R�)��3�]���]���a�o��M���.�p����݇����]�l�[�=qd��:�?��B{�6�W�v,����<�<YP����Y��T�=Ku��aelm~i�Cci'"]>I������J�7%ceR]~����m[�Bkׯú}��.�)'��v�M����ǷX狡$?��8�ˌV�Y��a��aP����#߉^���s"Kx$ʹ�?�A /���D��de�w�~���{��,�׊�b�\��6��}d�7�<�E@�.���賭k��eDw�=��p����3k|$���2H|Ջn����mloj���:@�p��j��Z{�k
S��fp;[ ��C`�o��\�3�� �|`*A�q"~���)I����������_��kf�^�R���@6�2h�g�.�%��Ɉ�_��.D$~�Y��>_c�\%��^TT闓�dǹ��'���6��[E�ɖ�����,���JY��3��)����b�Y�q�ΆЦg.�q��C�x1������_ǰ�/eƉ H��|W $%D"l;��q�����Msv����Z��I�M��
	v3}#���EC7ށeL�?ER�l��"�'·[a��HkU�.<3�g6Ϟ�6J<zH�M퓮�#���ް�e8��z>G[�k�jf�}te���!����n��&jV�K�_�~�,ܶ.ךZn��Υӡ��j)�޿�?���C#�&���ޘ�,˥�do�FNXRvI=UDV���)�<
�*0脆3A�'	Kv\F�����-Fd��i���v�o�l�۴���\_a�$��4���&pJ2A������=*R �4��g��l�j���'ى���Xb�84:��y�YГ��% pókƼ�9s�<b�kgn��8�(��x;�M�J,��6��8�Ҩ�_Txz/���>�.? V�q�(�������u�Оg L������m@�:K���*�0�#�m�Yy�`�;��"!d���;�B�?�G�T�Z+�3���9���D��!c��L9yM��'�w_a��w�+m�+Y�3�{����P{�/9���P��)��o�
-(2����¶6>�s�lB�o����^����/�	��_.,�T�)"��ʑ�I�7�Րӭ5�o)z�3�6$�/ɛt
�V�H�k�-E5F�RLWo
 �?����fj��SO&��lM�~���t�@��O=���0��m���X��la��2{�����2�XL8G?�*��2U���B�Ӻ�����V	�8�_s\��5^�Ι���3ۻK8[����"MM�l�_�`�~���O1���5�a�C0�N �.=������ـ%�oX�z;=��4�H� ��~\
�4�d��K�G�K��>8�V,��hݍ )�y�-��(\	<P��U;��#`]���V�?xU���7�ݲ�P�3Q�
?�!��#�l������"��R�uP���L�ǩePI�;��Y��(�2�l����:�L��=xp�][=��Q���� �6?�X�L�A��t�~<	71uy� �*��I�����h�c?��)�%�e���(�������b�����A+~�}�ܝ�R�k�W�AYYl���0�V�,7�!1k/��9q����F?����9���%t��"�w�X�����{r��f�t��1	�A����BŐ�h��(f����U)Le&��G�Ip+�Q7{�*�.�2��ɨ����Ύ��"-�>�G�#�`"�.�z�(��ca�Q���Ba-A�B��x�5t�Qp���$f�B�����y홫��C���%&8w]r��#�)�Ǎ��B
��e��F2@�֬k33w��C��O�1f�A���1}��$��(��BO�m���9�]�D,�#�<} ���
A ��}
i�� J�V��ӂ<��0�D��Q��1I$������,���S�{���j7L�wa��Et!�������ś��C��3����pZt��u>�Fa�o���Zi	*�<�x/g�.pؒԩ7ʖ�٘ڢ	��1ړ�\Q���}?0�@Q\M0-�JsT�?���r|��~Dw��g����MLφ]�R��q}��5{޸a	򇦓�P��5��u�윐�wERS(+'w��_A��	��0V=}��z\+ �F�V�)ֱ�����w��N���)Œ>����V�<�E������4�{�;�@���;#P!��Ш;.�F�	�����Rig�`b�nLA^��.�C����D6�Y~��ǳs�o��=�3:�׶lm��	��s�1C��:��Dz��&@�q)a�ݾ����aH�p�{t����Ώ��Ɣ��w+OJP����eP�ߤ���p��R��"�k\����)��-�p��2F��H�X��K�`�]�-���1�]6o�}F��O۷|�1Z߮b�'}��Q����`���n\���}H����E�9�T{ӝTnɂ�"�\E��6��`R���%<0��4�ހ舿�D�<w��5��)�S-��d�A�nm�~;j�|��_��5�!����P�lE'Q���{��g�W+��<p���⭫��P�ͩ�+P��b~���3�?䡢��VW�x�x���*�>���L�U>�J���G�3������ͳN
:!�Ͱl��G$ ��+.����H�����(�~�O[)�d#��-��n�b���B	��a�%-:t&�r�X�ѡ�P;�a�~�9ۭ���zu��d�9�G�)7rގu�;�;4���u������Fo�F������>��d�N1���'���4YPW���ƀ�LyRDe��vu�־x�����e���`��4D�wh��ќpۨ`��v�ڴ:��> �����7&���݋�k3�`j�Tx�� y9"��pv��\�9�J�f��d�U <��L�J~�E��}1u����u�z���ɚ��]ŃQ�_Xa	��~� 6�q�QD[Y'2r �'�*y�(������+�Y|\Y>��G��`8�ؕw��ӓ�|���1W�1��o�kV���t��^}#���x�&r�]��x�;P�,w�;f�R���ݹ�9F��������ZX��sŰ����)H7A|PC��h�����+�xYoijQ�T������fR��}�	�X[v�������\�,�|-)x~�]�~ꇴ{�׹�:�u���hW[�	�P?�0��MU��^ɹ.{�.BYD@S��..�N��M�*8��b�q-�)h\���0�DL�dӼ��:�<�ޘ �0t��]��p��+�HF�r���nN�tQ�wN&�#u��e��}���F �ծN�oE���oo� �����vrs�{��MR&.��&r'�*����K��R���X�7�rr�^Pu!�p��
<��U�((����RV�1�˰��}񝮆�~�Lgp��?�ޕ
��Q�V�Qߏ���ڛ��t�|�B(�q��:�O�A��	$�����0:E@\�1$T�#�.5�}�r���'8ݱ�P!XCu�X��Ȇy>R%+y�"֦$'�&�����J���۲M�װ�i���{c����#vo�XDVd{��a�tR�0*��]�3��2����+�i�M�.�Y���b�Z���Jʞb�$A���G��Mb���_nH~۰��6ui조A�s@XF��������:�V�@�"S��W�A������]y@���E�e�����{]�ј"Z�<�����7R�̪do����� +��b�fl��}_xC[K�E���(H�����}�5YD�� �q-eţV�v�#+�P���2���S�!5E4)f��ui����V(�<�< ߒ�2Kѐ�r�/���a�>�����Q�:�:t�5`�l�bH���D�����^]S���`�y��k8�F�(�b��?�(R�&|�
߀k�W)k)��5(��A�����=HX���ݴc�ܐ.�ٛ�v:��Қ�2C7�8�P�LQ�4xËe)�q+��S�[b!�!�[��SMLN�$��:�A`pō�/]c���|L�pK�3~��m�up�@3ޝ߸��H������~y3R�ˀ��jO�W�%��� �s+��]V+�P�5���ñE/S�#�Bn]f���
�F�'��8��"��O�u�����6ݠ��)��m�W��]����OdTZ&ת�y�-Sa�p� �DZ֩�-B��#����޴�M��g��/&�8�����2�D��yX��>����Qt�SE�?��0G��9��qNt��|�Z��D� K�����R<:��ڥ٫o���[߸O�~$�q�Cfk���(4��6�g)��2#V� � ?���T��_��<v��pIq�iꭳJW�N���q�ux�9��3ּʗs��J�Rc�×S�q^\����e~bE�k�Mu�8"���b��H,��:�~%?q�cf�exB�Us���}��ihyO�b�V��N��{�r���:6'!4CwUu�"Ѭ��K�{�A��/3M鷥ů��S|8���r���t���x��ӡt�&x��S����6g�k�t-��^�P�J�V>��W̤�]@y�#τ�Px��q����w�[�~�S�;�i��H��g7��;>��㡛W��������r���͒uA�o��v�M�g]w�2� .C� Z��_���v��������f�<���>� (U�\��y bu9��V3e9���$@K�?�9�+9<w�N���$=�mw�Bh����T�)8<�y�n2$��"�B��U�f�)B�����
�Q-���3g�]j%KtRw�F�����U7��p>��<2,l-��IbKHuIi雼����z�nS�k�R�TΎ��3�%���5������{$)w��s�_XV�u����;�O�U+�4�6�]�Q�|�Б��:�M�'�B��N|����[zU3�K
������� h�!�\vsN�����2\õ�, �/�����h��"�w<�:�Ҋ�ZM8�fRF^7��9�yα��uՕ�3}ʁ�%��c<��r�����v�(y�����丱	|p��	6�K2d�%kf���e�������C"xh��kOQ��m�ك��adN1�kD\�Q4�6FV�v$��aë����Mq���-�[�[�èU�Ba�
�M��h���ЂX ����B�Ao��TU�?K��,���{T�$����������s7����F�U��"�Ʃj��(+W��3�?Ҿl>Q��(�����*d��1�bh�^_7��.�E�OUl4�����1��I�E�s]��K/^���>|�F�d#)�A�k�My�M��:��|����z���TC;����,� xd�}���smGkh���a��J�K)*!�_�`"�˾�����>��?{�jS=�]f:Z�`�7���Ѥ����H5.������a-�G��Be-m����� 裪��]<)�d9�ԘpP�U��}�
��1�t^ȗ���&��M�zfvz�jh�_R�t��H�p;8�ɳ^w��yS��=j�p�;0(#zL=���\�2,c�ǔSd:�Pr�K�y��+)�r�^#~�m���Y.w��@�>"Q{��#p�~��(R�ܼ�lso�AB:�`[L���:��wn�Êy#�c��*��S�ݴ�^���l{H$�o�[��7�U4jdP۫��G���(_��)I���^��k�V���*��&2������7��ʳ���O]"e6a�q�lf[{ }sޜ�^v�DEC�ǫ1��vR�t�!6$�aޝ��1��L`׼�^�Zpћ�]�n3���뛎38Ղp��}����ޞ��盄�B�����Ls��"?b�3LP���jK�2��\1
C�񤄊��k�`���4A�q���x�F�i�*�P��
��S��5���8����e���1�����GiKO9��#q�����y"#Ư���e]v��C�mȨ"�#���R�f?�M�Dt��f"�0�C��a&8#�A^1�9mou�S���@OU������=GX
��ôu�SFǽ��uڪ�O6���$R�� ?�9�t�KLRL�L�=pr�r�V��x�n��e2{2��5��Ag���*m�'��i���Zɼ�-I��@`�����,�:�������M�������KWJ���:p l�(�w�^�p1�K]��iF�f��o���_�6r��p_$B��fk�5����eV|�)O�HZU2�>��/�A�c���0��^�z���&���N�n�!�U+����!�s�ė��sm>�S�S���A3�~��m�>�>�uRl����,t�w����BD!�g��9�^(�ݘ��op_�z�f��n�Td�3��?�X�g2�,tGA�7��B�V�����C<�W/�_h+̗��� �ym�9�
���c��k}{��6I�)�(��V�E4�Υ�3�ےu�.���v�P�����PeG�иX�
��wi?5�(���(����S�uK䱹ĝ�q���T�3�-K�L�V��=�*��������9�F�6���Od�:�@�&��(<�N�~�|���Й�<Z�,�44��3�Xs5l�ס+�#�7�����=H]�GT��Ł=�j~��rMb�>�i5�B+O5/f�q/*�l�x�!F.�+w9�Э6q�Tr��N�<���W�5�蔄�g�M>���c�]öa��|�V� ������'���]��2ʎ��!�Nwc��W-�����7��g�B��������h�f>dC�	��@"|g򂅄S:=5���oƞ#��,x��z+�x�b�I9��0��nm�\h������|��`�I����/�91@$a�r�S�����'ǝ�KUǄ�
�I+�#��k����
p�Yic�q�q�����&�׺�Hf^*0Q�\`$�v����LE����pL�V����埥?�He���:N���S�ԛ�03H�e\�TcR�
j�`�ǁ 9��$s�^�dԕ�����A5x�R�����a�����Є�=��f��li��$����T[|�ek\�!����ʖ*: 7#8���ۀX���8���C
�y`�ԙǝ��Ie�O6G�I�6JSG��+����gk�Θd$k�C�&�z�����͛���z;O� !��U�����V�V�d��o,�wL`��|�Gx�l�] ��<��2l=;cjum5&*����py�MQ)�񊂨U� >�&de�%��>���7���h�āU�ME"��°\I�@a$ᬇ�(7��	�6^1
M[#	�)�#u��/�օ�)4�K�����؈!ʳ��<+�a�p�L��*���3O���WCS�us�%�խ�/�sfiB��>�����H:S�N�w�*vQ�-��|��꠨��D+�3�	��(d,�r�4�C���b����\ߥ)������n�f�����EO���YV���}h5h8[����!��v�3e&!$"�A0�}q|��X���0��W��_�u��IN�Ul�?Ď8�#ؿ5�l���8���%t�F
��ck�e`A
	����bVV�
����[7>n�&�.q��t�Ex�3G����^U2�^�rE߃��Y���ēO��SoY����ع�r��1�磕�-v�`�@�����������}$	r[(Y^=9FqX�X���P>�M���1o͊G�?G��{k'���~��6�Oj�5��u\]zf�%)��}���y� ���9*�0hZ`TP̥r�L_k�?�"ӈ�Q%1i��a�u
� �D���0銿G���ue`8�)զ��+��ɵ܍
�z�II���g|m}:#�Ѣ��?� ha�L���Û7
{� ��˶��N�Q�� �,��m����$���M�~Vw޹�U�!���b��E���<8rZ�fs.��Ӄ���m��.0��)N}��<�m�����c�ɽ��M�!.�"E��ӿ%�nt��E�d(m�O��<�< ׮�{�u�*�»j�C�&e���V 4)f<��	��n_B�Lc��]�#��ʯl
�Е �y�MH���j��"���9��n|��Wݞ֎"d9�2n�r;�������k0\�;K)�@�\�E��&�?�cf��n7��G�&kӨ���zw����"Õ�7-�
M��j�C��C��VޟR�6�$�֣�0N��d�±�����u'a���O��$L���b24����u������V�D�H��G�=ӫ�X�x��Bn���I������xQׁI��Y��il�8q(�[A���Ʃ|��9�!�����L ��}�&���[�V�aH�uc���Ђ'tsHTݵ?g,�?�RI��߹ D_>n�1���S�E�������\G�X"���{\6�Q9�+:��� Y���&ɠ��tj �L��(�a2I��t��*���f� 3�)�N�}X�^,dͱ�r|]�`&��*L8,��l�=��`�T�P����,%�&���EP��j���(�4�@��R��U	���<:jG����Z�f��� J�w�(�+ۣ��ZB>,bOEk�p��vN헔�x��u`����	���#�ݢ~����Ý��y.�T���i����6�(����g\�PMu��O.K��.��k��a�t�ʥ�4���#YC{gǱ�&�������2�%�[d�f�qu��7E2��Z� �@�͛a~������.a��9��VC�.R)t��v^���?hJ�~�Z	.�p6��^�P)����Lt���O��K�`G����$�rK\��b[C��ĵ�2�Ŗ��K�tu�i%���Bg8Ws�����Ѭ]>g�A�Xs�6��(O��8�T>@�ӄ&!���UP;{&O��N�}M�J�8��fo���c9ȃ4 V������e��������$��y�A�Ǧ`��K��h��l����2dىn��Y��t��8 㻳}/�0�l��� /<`s%�Kf�CN�?׵- ��22�rw[ի���4�{X]z�^���y��0��l}��Ͻ&F��S>1����K�e��Hi�����Z�ף/� ���e��Y坫L!�ۥ;�[��U�/�[���pT���Т�_�;�Y8�����ǨV��R�,��:Y����@�?�[�eh�֪��[�������#�|�$����
S�;��a_"��aly ��sep
Ӄ@��2�%��3��IUE�!����v�_�v4z/Y��+��ֿO���Jz��A��H>�r�T�Y���1CB�鑸&w�j��̢}3�F����_<bkG�Pgj�O9%jޫ[�Ϯ�_��a���w'ά~�GM�N��`I
� gi6�05[3��!X�o =��z��,j��_m^�� �D:�����%��Mz�M+�^�m�4���Ηj�����{�rVb�챤l�B/1H�oR�ΑR��+m�����6a=�f
1f�г�V�]Һ�L�DY�KO���EF� ��Ӛ#Ko-�-4�����wo�9�⊝.�]G�O} �OnX��l���ŕT��D30$Zx��ƿ�e�O���c6]�al�dc�{2U�S�<mu�\`CQp=��՝�������a��j+ڵn�?3)�X�k��ooa�>�G?���d���p%Z�#�U����ٮ���J7,��§�3�R~$Yd���:$��sZ�����g�]#�y��kdh����M`�YՉ�% �a�[�w�Ǩ�G�|�J�?��5*<�^��� ur�㯒�٬[��7<�7^�o��3�Kh��.se�".D�����Zb��\9r��xJ,�l��;R�A̮�M��K�R�CI��&,�ǭ��K/��7�mE�"&ߪ�G��	j焑�_��,&��u�֟ڢP1A*�#��clH���}^�N�k�l`�W��\WM�y,#b4H1��F��x�� he�E_g��%}����J��<3�kry������@}ɷ�+ߥ#�"3c�NX��g�>s��:Wr�J����-`���>���6�����L���l����s�߭�O?Y�P��M�wR=[u�,v��b��5C�UH4�~BTv��O����a����Ol"�o2�}u�{3�:�ɍ�+k���6N�q���9�����O��bf���8D>�)��?[�ޠ����U����|EoJuj8_/@���$�~�t�fؒ*i&���K���)ˆ�k45�NB�_��T���U;�s�͍��]�.D!�}�.'�-kW�$ �-g��P壦���B� �.��F�z�ϊ�A���<�W0�4� ����B��Y�u���,z�����i��pߚ���Ē6*�>s�X46�8�]�bB/IM/(3�>C�4=���ȸ��P��Mq���+UiXu]:��Iv�ѣ��/�*IV>T��=Փ�k_9F�H*�k.��/M>��-����������	]@m��g78)�-��RZ�nK��'���h�fK��&�!���}��\�슋���G�ê�����;ދ�Wh� ��C�Fs7�~.�>���fm����%�`'|�l5s�Ӈ���B��P�y
��C��>@����@�$��4�9G���%IzFrwZ��J�5�S�0��Cj�.k�B`��ǷREr�ԫ��y����)/' ���"BqظP�H9	8W�C!�@�S<PB&��d�=.�����z�'	.��'�+=ۑ�ex��@��r�H�\F�ي��gC��>H����Vd��)�����@���������֓~e|��v�ט�C,����}��5�fx٘[����h�`�*	C��N��n��#�������$�x���e�j�Ƴ�G{U�[¡ӀP�o t!a	'��l�I&?U+-�V'��V�t�ӥYP�\������2�g�7R���$��F�n~��������t~r )�p�b��yT�-q'�D��p�NV�0f�T���������"C(%~�~i6p��q�\�	��6��o����{@�O�΂�:q�U}��Q�������(�V�Ē�� �r �/��a�ʶ�>�̏kQH����V{�ea�5�;:*�5hg�M:I��DG":vS�����>~�	Y��0�]DT��NaY��2Ƿ�ւ�٥�?m/�
�m@SZͮ��ʘI��?���xs�	Sw�h�F�+���g�ؗtg~�(�[og�����.��Tם��0�|ȠUza�WZ�|�`N��W�j��#�RJ�곙�9�B<_h���M��5]���k& ��p�0��}|j�M;��|Zei{��
��LM~=��vsD�m)�W�I��pg������C@�Og���)K�� ��NޯUg�xGh;"G7y��3�d�X�ٚ!�NҴE����o�Uom:�祐J��k�'�����`_��i$W]�[I���R��;��?� � 3�I����n��(
	*%����bs�����!ί��2�5�~��M`��I��ꞝh��{���C���g>$:{����������'��׿lY�Ni}��O���3bq��6/ɶ��:�!XLtC�o��r��qg��݆�O���J.�|�B���-�P<K9�R�� �%�'�M�;!���<q��_Ieip�V5%��>��[�HJ�?c&j�<,c�ʻY]����&,�ĩӻAc���K����}1����?��h�_����=�׍��Lp�����4�Ђi���� �Y�]��F��i����~a������D��Ɏчt�y��H�h>
2Y�{J!�9�dה����ҎN���d��Ǽ ���Μ� nͩ���e���`|ֽ��V�?�O�o�<�'f�z*d�܇ZDv��c��d��')?%8i�B+ј�F���U�c���@�O�����=�;�=(L�ň~�ߤ��0��Ճ�S�&�:�9��¼S[��|���wj�
~ت.�V R�ʌ��	�; s�x%�U�+u^=H8G��v��E�Ǵ��SB��{��)�f�����KL!�Mq]:�����g]��T?��?k�_�ZH/*�r̐�q��
�W���N��(k���0F��vد��zR(�ϩY;+U5n��2�Y�1����eS�����q4{����
{��
q�E��;�����x1/%�#+gȍ#w�_D�sJO�hsi	��`�}V̺�Vs�e�5M�Ї��8Eץ��3vNB���gj��4������h,�늘JY>���p�t��\��QZ� l���Jh����e��	v�ʕZ�~MkHS(i��N$E�����M]�#_��HA��bd~t6g����p ��Mn���e��#��'(O�&�J����f\Ƃ+]��!�q�m� `2��v��C��_�2��c������5ܥ��y���鰃p�s��ѐ�n��i�+��uA�TNL�>#73��[AH�EI2Kzv���`�gmd=a�(�����{&[hk��*���~�/g��:�6y���jK����2-���3?�P+;_)ַm����ā�ۑw�~���]�H�]�<"����zB�V�Mh������*�rn$1 ԙ�I�>յ9A����]�! #�������<J f��O�ʳF��Ӵ��L]R���e x|��lւ��R����nі�z!̇nř��$7�1)<r���`&^QVE�yL����u�a��<Ij�*�ޭ�/�b���M_=h��už��۟�&����}h�lP�1���3X�C�3����x���)���o����j�cX��-f&!)�u;�Oڹ5b�x0 N�L��ܑuj��uk����l����^G�VD�\�zxAA���?���d�N�ng�Z�%ܚ���98�]e[����$�竅<��8���;(�"��6�'��=_���jĦ��� �/-��K�{6��3�׈b����')��v���t��?w�Y��A�0�zn#��@���V(�������\�y]	�(,�-�c�x7UvKȠ��"Ն�/^�E+�m �
a�MX��,3�s�hU�F���]}�i����!�Q�(��d�h��W�$&r-Ļu!�� "�&9����b���@��t)�[l7�S͂����h�5Y�G�j}-���`b�:5�>S����b��g{��_�Vd�΃��i^�>�4�>��\
I�O:F�=_�>tb����l�Զ�s�i,B�L���r�(+�;g629H�ah�v�x�"d:9G	���p�_��sax�>�ET+[#���T��B�S<r>ȝi�%-R�*���]EI:JJ�In9�W�D^V�OO2#�D�pY�nR+W�l���K��ꛃ$���)��A1�W�+����)?��ʚ��w����
�ķO[X��1���4!��-GUOVǋqh�&�X��)ti^"DtK`� y$Ϫ�4j���B�a+\���Y��c�cF�j�����뾅���45�Jt�^�7��Wnz�����x���� ���M��
��y��x���4hR�Ĺ�o	��yq���2a[�0F/V+E��K�餄� ����&ʞ7���X�ow�Q����2�>��)�Gai�A��)����,�u˨+{:����Ǭ��)��',���!��1Y��fЖj�}���,b�g��3�ڃ��H\��>����
ɺ<���L�q4���14V��n��s��7��������'��&�Hݘ.G�O�R��1J���כD�^(1W��ظ���׵R�	̈́�^�/5+0�B~FfcFF����[��&L+�+�ð�1�g"���$m�` )�_=Q�{=�ͫ%N�$�j�=���DsdS��K��<'r���כGk��CRv*Vl��Lv]{����P�E���)�uֱH�1�����M7[B4���S�&	c�{D=_jD���p��s:�A���Kjҕ�7��l�>$1�V�&4��޶F)x�_����F�5�pkҙ�e9�p� ��8A��asF4���f��D�S	q̺�����Ht��)7����U6qq_E�3��(�G�Kj:d��.����U�l7V�b�b�f��$R��|�s`�%�'�\���Ћ�g"�0�qc�ҧ�Q��oo*���cX��i��\I�|z��|����"н��ґ:�P��,��e�t��.�U�aIb�G�Jʸ�C�� �h!?��)��9����3��f>/��}H8	�̩{�nH��<J��Ou9]y+l�u���Z\���_T:�D� �O��4�&�Y7Mn�Ot���������z��9�D#�����e*h������P�t�^&Q��Q���XD�x�5��M�"�=D_��V�Ɵ�v�&�f��p��dˁ>'���~Ӕ�n�eţE��͒�f�)�`^��"�:2\S!|\��L�Ћ���l�d��6��(d�g�⃕�� i��w�+�W갖�WO��w�eO,��y�qe��=�m����|*�c!�2�% g�HV��A��!	}x����Ʈ�}<�Y� )^�G��-<z�I�4z���<]bs��p���.�¾���h�h�rdѝ�v�ѩ9��g�cP;ԥiQL��&N�<�M�j
g׼���������ͰD3��7X n6;�~%���<�uL��g>��)���B9������GTO\a\�B��~'��kS�n�����u�>w��>���M�E�'o
��B�<�1�'Y�zJm��#����?(͔U�;A��G�̢t~O��R-��k\���s _v��ѓ�Pc�g�,����cKGoV��G�YS���i'�O+is��*i�E-�Op���#��|�7����)��2�h�\ c���x��M+!i18�Zʰ�}�祚ԟ���))NЈ1������8���w�E���񥠾NݳͣQhf�}L�%A�p�۶��'V�Q����|�Z��HPMʈ�?Xk(�|��]-N��nqak\,�nQ��]�N�� !��N�����_H&#@d��~��[�3�sK�$+99�"�����;�"/c����*�۔L����m�i���~�����k�:��f\� ��}�r�����#�R�I,�>�U�VSq`H�E�� ��M�u) �Dfɐ��N�trh�=.�p���_a��=�(���L/����V�@3C11"�z����vzm��T�'��-z�I�s��������^
��y<U%���q��7hY_`_����;��D���?�G�G�})�s�
Y������'6{�֠6�e��U���S�@��&�ai������?M�I#������9�9`�t"��dHq�� ҽ�sm�F���/��օCP�Q�����UJ\H��	�@7r����ힸ��=�0`|3�+.��]d���i�8�gьY<��V:�7l��O,��N{!K;b��qM���tth�Y5�Y�DY v��,��cf#��C�z	K{�m��`C�[�4��kh�&��j����'����~
x��[������F�9���c�H�ү�D;�)��M�G�M�R�=�RF��z��"[��e���4)�R���/�Ճ)л]Z�|V���1��� �+SS+'Mĉ��3�*��A�!���3��jp���(E.�j+8�ڸ 2�=���'�^��2�lIA��d�l��4h�6�<�^�75���������m��ʬ�H�X�ZKQ%�V\&%����I����i����Dq�8�wc�`Jq�;�}.-�U�~�Pu0�Q>F��]Ш>�V����
��*�+������Щ�J9p!�W*�̠0CF��*�B,��_���x�T�}���]��=�{K��h;MF�.MԷq��&v._O��D��=�*!��{�ʗԥy�C����@�\L��.���`�{3"m��*%N�{��|��#��Df���i{�x:��}���"�!��&����*�4߿������Lx�fzMrnx�>�^�U-EI�O���7s�	L}f��n?C~���Zj�
����o"T0�(���L��FI����Ŕ�K%�"\6\�]�/?��'#�8�e�L�EB�4����'�"��u�<Dj	�_wK�[�K��@xi�fҺ���;�
�HT�}�`O`.0OY��z�i@�Q�L����I8B�K��ik�G��;F��;Th-�p �<z�N���3I�!��`�;!�]^d�|NU9TwF�؍O�L��z�P�ze�gg�J��_��W��'�3D��Z�FG{ 5��˾q����x�0������.�Nx�«b��:�r�1���0���3�k�<P���S�C�����釧շ90waE`WҺ�G\��?��E�$��@͔ f^��8���l_c��%�=1������V�-�o+Q�V�}G@����zLCD�_��(�r��,_�䔍l����Ce�<�"����D#27�j3
��̯zS��7�BG+%wΕ���"��t˳-n�U��V���'�+�ӡ���4� �����7[��ۏ�EDC&����q�ֶ�����X͋����eg[��җF�� ���&Y��1���R�Na��$X�.�b�Qi��O����g�VN��l�ik�(��8��{����	��4q���0���
w]��y)�����۵���&�<�|�lv�3=Zf�c��f�=� �Pމ��֪E����`Kީ"X;��#e�����Sr~�aV��d��T�]�)ۥ'/v�����Z��`P�**�>D�.�ƾΌ�ķ�����M���<=���d��G�ii,r�4���Ǽ�u2�p{V�D ��kH��3�T�~�	E��m`]W�ٟu��aCr(��.��s���x-��g�{�J*m7$��Ca��9|�8�5��y氠'g����g�	�#&���J�İA��׆2G���F����?����=Yĝ��ݿ�ｖ�����$[B�d���E�X:����YIy�+8.ۮZ�|�Ya4�KD�?�~(�~����!X����1�Q�;6��5s�-��챲"�:�Zˁ���9��J�Ǆ�	�y�Vu��%r�F�?�vI*w�"��7 ���}	�^�Ս/k�|M4���s�V;�%�\"\{��b�r� �ؠZ6�p��=��,U�Y�5FJ}az�F�}M�-�f.N�I+�[ ��Y؍����D8q����dY�"V��_M"Ġ���y��U.wHI��}��\�14�l�j2�I��2|�?U^�Fx����%/����Q�g�x7�����`����ёG��p���@�h�T���t�Gl�'�e��tm0�#���w6�-�_6�Z$�P4����r����uUHW6�~���%�'��ln�X?����@i��� �IK�6���#x�<��@��nG'+M�8��D��~A	0U{Qe6�b���}0�|١�N��|��=��U��s��J��@�O�3��0���^�N�� ���X�ě<�XŌ�
 }/�7�~�
^�{�)6�v�����P���G)�H���W�f{^dAV
�Er��at=�S��+�CO���
�O�LT�DYn��"�.��(m���W�� W���' �8�w&M��$x����b�_O�6�y����E���`��m0�Z
g�,�:��^M�T ��5=:`���]�)����{]H@ �1%Xv{�����R+�X��a�g*n���w �=�|��ND���4"�d�=sN��wׂ%�0��T���B��!5�A��R��kũt>p�^FE{0��隆ol��ؠNM9��?ҙ�������Qnҧ�/��-[�G Eُ��{1�� �I�>�#����C�fӀP�����b���ȣE::I��/
W��Ȑ�E�#��^𨳌�Ɔc�ρ~�������H��u��P�L��[4� ���4��%_Q��l�\�+�&@O��6�I#2��+�p�.F=��ֹ�k�-8k�CRlV� Ed�d�0g+L�r�
K��p~��!"y��9��@v�h��W��lj�9�r��Ŧ�1��I��۔D�Z8�������*��	�"�6���_ v]�P�Y΀Q�����^�?�y"3�Z����&R(���v�a]l���&�x���J&����o���Wu���y�Hc�����/�e���K��Q2�`K3�� �uۂd% ��^7�\�1�ۄX�jnS#.�%֊l'K��2�/��Kq�ς�ܣ�.s�OX>���z&�m=K��R��j�'j�&�᐀���W���s�P�^d��Ϛ+p�B�J'P3����B���s>���yח#���P�!(	wړw��TN��e���^Ǎ��;=�P�P`BEr��Q���/��ۺ'B��$,��u����\$�'�1�H��'V �BA4i����_�
���	�f��F����t��-\�%%4�e��lh���	�*%��l��Ҡ�,>�<��푈�$�R�,���\��@�9a�Y_����0��ᨩ�,�"쟑�܍~�����yy��4j��9��P���u��{�B�����eC������S��L%�f�̊��x��>d����u֎�E��a�ty��[�N�eZF)c�46cq�QAt6L���Vѵ�,��� Dz)��J �@ٝ��m�wl���c�
+?�m�P��&�!:���a ��ĳݜ�t�Q�U�ڽ�q����amA���������c^�a7�<�9;U���wPЅÀ�o�T�~��"���C�����ƀw�!��v���M�����/ E��a)+XS�@?���z^v)��G6�P~/G�"c�d��������52�f�v?�rwN���;��͊exH�W5�YOT�d�b��2�*�������Ց��$b�j�	cwG3JE`.�C�SbO�w�5ƾ#��6x2�x`o�������M�0l�g�ni}����тn�Zg��0��S�e1�=�"�9t$�m����u��7��c�i4�4u���p,4$]�Z�Wi^]�i̔����"S���$��DF#�Oo�U��7\�G� ��;��e��_�%5�y�;©���]lA�	8X�2�Ē:š��v�-b��๋��k�p��<�'��o���"�c�+q�m�Қa�2�&�?�!��ql���H���Ȧ��2������}n���QPԣ�f.5g�%�&}����d�g8��cB[�!��� �ɰ&J������0G��r�IAii��̈́�C�Zh��%
�
���I�곶Z�q���jiO@}G�
;�s�4���r�.�5\����l�ճRo㇄\�h��� f��1�=�D�$ !�ђͣ�g�/��t�������5�ݭ	�����р-��=M�F����<����G�>u�	�����rsx>j���U�˒�p�S�/�4[�Ź��n�3�"�K=ʃ�9�I�F�RI���k�H`��'4�sP�Wf���BGj#l1�riO7�q��W�!�G���8^�z�l=��.p]ņl���7��I�\�|�82��r7$�v�H�����+���w<�Ly�L2��sl�&���$v�)��{�G&�#�B���>��k\�@<�kj-����x3זq�k�ZJ�eG��p�h��B�E;��>h���7ˤݖ�w�����fX����-h�&!�w�3\K�����R�f��yp(����
H�$/�6�r����^��h��D&�����=R��9���;�E���Ճ�܁Rf����|l���/1���Os�?����VC��JC�C�9|��U�̈�H�O��b��b$����=�2aCg�8�-<��9����r��"_���S>�W-b:�Ƨ� �����;��ҟ_�b��ig�{;?ȉ������ļ����l'H¬�u{mCOA+�0E����h�Ðlt�)
.�X�z�%��]?ʅ���������C���޴���v�n���a﫣�D�!&��c�6z�$��}��ً��ǻ[�t��� %u9���~��&�$W�d`ɸO�!�<ct �5N%N���Z��"P1309�d%�H����m�]~�"��G�[��+�G`���	�QhB�zc�oMJ����Vs��^#�n��}��rJ��qs�A�Z��j�1eI.�Y:�Ԃd�U���h�f�5`��(��tD-@A��M=�^A�i�{%��;T6J`mg�(����a��I����Ԑ�!�\(GFVG��Ԫ�=3�o��D�D �c��J� T�Ekt,����T����y]��2r�D�(<.�D"�6:����h�j�k�i'B��TKg�1�
�O#G�JxZy�ҽ�x�a ���ŧ:ς�:�䰠����0���J^�8��ξh���g��f��e����	=w]��QT���X&���t��uH���a��=w�l+2n�Ԇq'�Y��;e�� Z) �I�/��̲�°��Y��';򽻞9�(�DM��R�s�Ш��r�,��?�y!.�j��#-o����1���e��]����I�~`b�D܆z�[���a���&l�-�Sw���͜��L� �ǡ�C�y-xgrN�"����ޫ�=��yWR����Ta����[^زJ둪���c��jG+u�R���I�kt@	:u�.[��?�=Xئ=��=�U2Ҏ��vt�@>	�.�MNFN,��H�^�G�I]�{9R�V�0+��5��E�I8�q&��4c��E�\+k�^fنXpW�$� J��&Z�s���/3�-���%��%�]2i_"�T���W%$^�ӴD�o���V8j3r�i~ӕ�[�f��̿��V}���t������#N���R���n���寋NaNW���aH4�yV@%���Y�;z4�[����j����� ����7�����D���j/�`�]�[�m�Zu)�-�L���Y�Dk�,�b�{1���?z����P�����D����j��;��S�sD���%��^�w:Pg���L���(8]+���� �5�Z$&�\5��ht�ZziR���r�+��(3�1�,@�mkE��T�ENdN+6�!��fO��.��y�m���w]��;j+�'�xpA���uPYMq���'"�g��V������mK��Ï�{)�VV�H�Z��__����4U+���\.�(�AUq�`ӫ���z弝��\٭�0-�t}�)��5�}^�]� ���h�5�SS9�iA�i�7��ۈ2纔N�4�����3�,Z>�E5�Q�xҘ�f��W�p|�12��ݿt��r�W��)
{�� X�|���o��l�.��F�?S�wc_J;�����-u�Ī��1�Ϲ/�ٖC��35hY0}��u�Ɲ�!tJ��(Űf�ėO��L��92���c���Z��O��.e�~ѩG	����N��dk�����ŝ8=���njH�Hx��f@�*"�D�������~�q9$W��1i7�u�)/�g��a4~q�{H�D�c�>Z� ��!�����B;��/F��}s�\��Q��	t��� F�a�H��'�ٞ}�R����5ݐn*!8;3�$#˗{���ɠ��[V'�@��ۗ�/]��C
���x�Qz���Pr+�̧�%
��=�nl���^��.Ƣ)7��+����
I���[?��L _؉5x��l�g�5W0�x	�]❐��u_�sش�n�]���D_�Z�J#.��7G-�yT��q{���-m=��䵁����!��IEx�΂�ZU�Y�q3�W��
�u��i����^�~�-�Mz�%�M�2��?���3��ō��jzҝ����s%��ԃ񞘸ko>� ]�� ��2�:�dB��My�������95d���䭈�k� v�]����3���}����ܽ?����5�$���mK>�}�'�� )�~���`�s�3��&b^ A�*��T��0&��\5�~����L��E�͔�ElUuiWu�Ǐ��Ed� R?���ȇ��4KKo1Am�
�a���z����N�� �dp�8�%�K��n�S��X�*�ȫ{$аg�`�VLg���7�#k�C`<�fBG*w����4</��3���<� �x��\�+j�
�/݈8]pU����05�1	i�J#H �/�]y0�%μ�z��/�w_�n`�p�RQg���}����-��˦#`�5!����i����^�%�z�3��✠>LH.�<7��6lD�Y��mЁ��rY��`�s����M�p_a��/sT��+W3,F�ߗY�$2�d��m+\ լ�B/�.���(�>;\��A?�vܨ׵��X!�9�~G)�9�ѕ��c;*�'���Z W��9���΢�&���+<�3�ٟ�Ǥv?�֭qtXTD}���u�ӟ��k�����N4��n�閭�$��n<�2
��3��jex���)�+����ԭ�#Lڠ�����64�~$R_ȱ�t�^@i�g�Rz_6}��āNP.5�so�	y}�ؕ�z_��$�^�wy�36�}��!�Bm@
H����-�����Q��0��-�n��g���z���AI��S{1�5�;ӑ�֌���ӆn`Ad�i���"� D�K�m�h����#0�+J������c}�n�sFQ#D�G�P�n�)�O>ɌI|e����%��O9���"�
Q[��
���2�2�'M�&�i���ahY����-��f�W��T�/����pTBU�B./�[�ʸ� x4ySER��Z�I�������_v����bo��$�P�:��0�����7a?�,��!&�LJ��C1��Կ	1�I^�S�O�Y:�Pe3��&L������z�tW�v�[��n���	�^XO��f�|�Gd�Itc=U�@^A����؀O��P�|��R~ZD�����9�2zəՄ��%,�!��>��7JÔM��7a��L\6$R�Ō���2��{K�C��D�QU��AlWrx�<�v%��P٪���c�-���k$I�|�?@��.?�ez��fܯ�/���N���~����pL{a��a�!*9[i7��;RWG��d�I�xS�L�TJ豄�8v}:FO�o���G���ef�K\x���~���KdH�CZ ���G8�u�9��s�>�׉�])ǤfF�n^�c����c�wFD�,&�E�5WR�q��#O�m�Ν��.�]B�Q��B�ۿ=P2�7ZQ�n1�x�..�N-�-�J��,�_��14��Æ�b8�*;%����n+�~�YM��>�� ��i���/�Z�/��tK�_���[����vC��_�F���"�jP��1�L���{e��bu��_�"�^TS�u��nn&(�q9(����,�:'#���2�|�!����xɌ4~s��sq6��!��Wz�h�@Z�ȑm����S]��H���]�߳I˂)i�9p�'Y�M� ��Nja_od3؍��g��� >�
|̭9�#�I��yi��(�Q�h�t�߄|U2�K��H ^Q����:T�su۸H�*���#H7��n��N�8��N�ƂIڱ�!:T�үo��uk�$�y��äd�U6{���'�6�勚 �j�5����:H�hs�ev>�2&�� M�dګ�t�˻�+��|�AP��x	����QY�j�9c,�����OxC#�l!χEgBM�Ԕ3��E�΄�e�j$|	�vpp<��īx��#�"9�.t�7�＠"\y���d�YV��P���՘P�G�Ija�|ET_I���fēs��Һ����9�z-.9�sF�2ĬB0��XJ#s	?-Hdש7�ۈ~z�=��J�!g�/X(nA�c>;po5>���E�7t?h<$6�����㫙S�	���C�!v���S�����i��gĸ�li_����ܾ��V��`�tr�ڝ .�&T[�t�`��3�`F?������/�3�/J����.dLJ��xQ2�v?�xcr���T����±l���0L���SZ6I /�GYJ��=d�iH��p��_}"�C@�{�)<����{y���B�/�y��ڎV���K�jE`b����>~���D������S�t�)��5Ҁ�h^��5�[��ҍ��􁪆���R�z�X�� �.���Q��q�q � `bc�v{�|�DY\)?�d��?�]wBd�QD��$B��ɹ��k��u~�%�H����\$-��.W]����Ò�
OQ�H��Eǻ�*3��7�ܶ��_�����s��6�����"�"[����UK3�5J��W{�z\6$���̀��oC4���=_'��&�]G�"�Py�'fo^�|�ko��5�� �X"h�e���ܯ����	�D���A��=墿����eh�T��Ԃe4v��xs�Ky4ܐ	)�����/��l>

jb�V�0Z7���J�)H���u
�P�jn۳8ջ݇
�p�?���R3\����)��o�o?KQ�'Bio����P^��c$�	U'lb#��!Hҏ�������e���/��|R�
�?DP�9Ju�����2��	�������5��{�"ٸ��6���\j'K�UD�}>yIz@����B_�eF,��*���>7��t�Q��R���n���8		A+(ړ]+}(���-M��=�A)��o�ݯ?|�Ι���"x!��ŕ/����R$��3J_���}0<���[�K-M;p���p��m��Я.�CPE�ɹ1�[s�����ĜjME�5���;���O���8��e��𧃇o�J9��ϯï|4�]�-��w��mEᇓ�;�&��dS&�"#3��R�����9ɹt�rIL�%�>m~����N!�y���B~�x�(���ǌ@.Y�2�����jK���}�(�����mdy��F;����~{Q*� �E��6D^48�R������ކ-(]���'cV1��G���CTs�5 ����&z�����W&�g��`|P�l<'a�02�_�ْ 9gAym��ǧ�M�j�T�*�
�9T6��4�l:>�s��v4� o�;3�)C�Nx���G�V�b&iKYm��b8����~�Ζe<���B�W���cZs��=��_"�Gc��ޣ*�Y��p��e�zI5����Ju�r%i~�z�����g��(J�(,��%W��I��i˃��Dru�q��y�hXV�٬j,�^�@T�3�N]yF-d�����#��MH��;���T�^�A<4R7�Y(L8����pe����ز������+�3��r!��C��ӳ������F>�ix
�Jח�B ���h����*4�@��]T�I�&^�]$:W`P]��s��K-����Z���ˊ�V-�ݏ��B�U�5��4?�jJ��9 �E'���xΧ�bL�+5�Vm�O�H.�ُץ�f��  AX���T� 1�5�.�ࣔ�M-�W!�i�o��<F��bg� �Z�bHf���!��￟��N������K�@@�~��\2[���3E�^naOo�k2֟��	�}�A�v��/7��e"ڽ��ıb��5ˤ�ɗ�X�w����u��,6�|W��UI�07U�D�6Nx��2��xB3�*����搭M����ka�� kc���N��u���s�C6��y��NK�n5L�P����,�3�@�s|�w��k��H��V��yv�R��z���M���d�G&d��"Hw'�#F �"�.��~���I��S�����W�׃)��K�5li$��f����Y�|~W�#Q�Їíyc�Up��Մҫk���[><۷@��0-���2鄘db����U,�����nc�*��:+�a�a�T��"5��~�D�2r=�WF������.A�A��e*Fj��
I�����>cm�����a�0k�Nd���L߈�Nx� ����{}�M�ߝ�G�ƵK�8;Y�^���M�����(�4����cO�|#uӡk�]�՚D\r����1&V�k��7#���keh�W��*x����4�����Q3x�Y>tji_`[���,�`��h��~�8b�XW8�9�� |M7t�������cձm�4�{<��� ��z����1���lu��!�*�x�s~�i�/�$s�I�LD^��~��h��`"SB�ʒ�,&6��A��	5j�xH%#��|�HY�2������c�3clm<Q�N(��������Y[�<�68�Qu^P�>hF0���I�n$��(�F_n��_ ����2�7Y鞮��vqr�P��F�P�G�,pp�O�e0/E�r�>�\��8�����.z34
����َ])7fۇ�&��%K��S���Q���C����+���}���F�q��|]� ӳ;�}ڈ�O�	��IN�`n�Avs\en-��Z�������2kc�G�t�N�<�#��&�`��\U��;ܪ.�f߶N�!ٗ�eH�x�@�I��0A��sG��zg��qo�G������
 �$^E��S K�r~�R��ס�~�8�6���(jO���1�1֬����E۰��/�W�����U��t)���} ��T�q�B�u�&��-��)(��cᗫ�|��Hݽ}�vAdD����$P�Dmu"�6��Y<�����Fq�uT�m�K���,�x��9W�=�x��c���X�s�o�A��=h[��"�;S>a��
K�)�xlP ݰta�%a������_|Ighr�%9T0�H�M��E�A��GQz4��P�g�S�%p�:9Pڮm<C K�`M�T�k���y3�(��A��e6
�ڥ��ס�F��tע�W�۞�s���_R�Rs���m���/�m��=])�,E�������5��S���b���}ŧ�KY�_l҈!;���〈c���2{���j���C�Ug�f=�gX�_|x�Z��d�L������fZ�L( %��̌��Q�#� B<�Fc}��^���S�M��u6�,����%Q s��_�6cY�j�2���B������gC��X
��	�L��%���\�Ƀ	~L�"r-$�B�ڝi�I�+�%{C�ѝX2�_�k�}{�0��a�^��qa��W�\Ю��l:�� �	��B+�35zitQӓQ�}Ѿíy�D�0��=L˴_BҾ�_�~��>F��C�D��V��6i䪊	�׿�ĝMU�� �`xL�n���b�z�,��O�(t�����'6'�TU�_]��ތ���jG�{k�~�C�{�	E��Y�8�`�836�L՚�[�I.?A %���6�-tN�[:�co�����=9F���g�n�� r
\@9�V.�yulAׄ)��
������{�d(�Ȼ���YP�(G��l�U"�n(�[pM��2���{�B���¸U &�Ѩ�,�\��9=k�	ץ7%�Ƞ�����������"���&��D�f�ԾP��s:��t�A�����ЙaZO;@��s7�YS�<@�K,�,���G��11m@k��D5�������L��Qi����$CV�#���y>��L�!v�mN~ ���K���0��a�l��H��������ƚ���#@���UH�B�Zvv ߵE^�z6���+5=��*'���Crm� �j-l;�k9q9H�Q�b_8�qL���� �����cS����>�'�H��Wy�&�H�;$>�)��?y�p=�ä������"��P�>L�X������Q�f����;�����#?�E�u^C���{w��E�,����3V^u��m����Nל���!w��d{\�Pn��:VL�ı?���3�H����t��$�ƴ�sD�F�����t0	L+��&CJ0��]?,��zT���qA�u���WzZ!�g�oh娌��(�������uy�.�8�ۄ�d����GS"?dZ�߂U\�ݴ.z�\%���L�0K�`����|�
��=�wb�-�}���
�uD\Z�tpJ��dT4�:�N�:c�����kg��DK	�A\�#���E�m�{+����j4����H2H��$Rl��`����n��Z����me��t�]�rҨ��ΰ��������@P���>9��z?Q�sJ������P�c��%�46����ÌA�@d�ryM�3� On(Ƙ��@)�T$���Ka�&g�
qOF�M�[�}�ܟ��
bwĸ��zU���P�Ւ�XC�E^�>�W����Q��5/tVj�e��I��߶oun�K�8������;M�43�	$�?k~��f����=b�v#��pzMв&8j2:��� �W���B.ɴb� �N��?�?�W��ӏ��%1������{KqyT�'F�b���d���Dtb9�f�V��w��0�0�%�5P��ǯ���c�;���C����.���)���Ȯ4��n�5�sw���0��Jf��{����㠾��N�#����<@�fѩ�R?�O�A�:l<L���B�z��;UW�#?s�<��e��'��wI�+�;�ꉆ�y�-��� ��Q�^�C�i2i$���C��6�ߑ�[>0" n���lX�&�!R�^���"����|D��B2��L{���*�ݙ��ذ�\� ��n�\���c_�#��!Zv���B-bx�?�uPF�B-������2ո�������J��c�GA�E���'`�
��'�����F���62q{��:�{8�����5�ZB���Ҷ
��P>�E$���|zDM�2���iV�_#�
�n����Hs��@"jh�Rpɥ�\ew���1�)�ŝ��݂{�z\N�E�xp��&f8�4�W;`9f���Hw*?��zs�G�L'EԖ"���<���:�0��6�6?<-Hc����J�c��������8+Q)�$4>O�������E�"���0��dTkUˤfO��ϙm�˷�q�`4 ���͒�j?Py(`�Wث��&[2��wl����4����֖wv�YYʱ֠K��{�onXw�f���`/���g-� D�}�f\}��0��6�����}�#�L5�)K~�^�ݘ�������I�"B4M��,�Ի�{&"�E�IIB�q�׿�f^�
���8��)suJ�4��am���'�l�+�r�ҭ�0�Lo؃�";K����T������������tcL"j�b��v�k6��k���"�ܔ@��v�Zw�r^�P�Z��~�F'�-��j|��Ƚ����6\'Q� �L1�DDlp�3�1�N����(W̚�o�[F^�\���_.Lu-xdk����a�k�kCEv� �y�5դg��Y�4yD�
�>��A+�)��z���n�8��M�r���ƽ�;:�����>�F<��,X=}�S��(�H�q�zZ�o�;p�2:5/.9wG�ƤPU)�o�'s}q�5�Ѭ�L���wؐ�-�fe���M����-�JN�
�b9:.C�P[�il��:-�`l�(#�@jC�&߲�����5b�V&�v���[Ƌ�-���Ջü1��Rz�r ����Sɇ���euF��AP��%�E�z�;ti�+z+���3%�]���5x���;�(�Sv�wq|�#N�.��ih��E#Vzv%��#۱b��Ј��@E�;�z5_�����M̏�a;�p�8�SKh�˯���7��h�/�C�V��
{҄��0p/7����`��q)�/�)�	n�L�@�Y��r܅��˫JG���]�q>y�*&��*1�U;뭻&VVn���M��z�p��6%�ǣ�ܻ�'-�fk�K�)�3�D��rs#�WQb�~��?����a�{Kv-_r�Ly�Up�SJ�s���9SM�'m܃�i>�:�`:O��J�;��g�|�&���އ�u�DVVhj��0��w���f�h��.���f�â�|١��G\.݆��xF�F�����u��SPw�s�3��Og� �̷�S��H��s67��[��$V��	/aK��2��A~����(���*�]���)�^,��]��$4^S��B�
�;� 49���k�(?������^�E�|@���!J[)�}5mIv]��U-�K�_-�%GI�,˔c�D]/i>�+-�'��+^$�D*q��
=��C��$����U��׫x��R��0M� I��A��ʶ��dɦ�=��m��x5?��Q�Nؠ�:�P͡ �C���cV"�	��u���#@��c���ir�'�jsv`��E��b(�	~r�� "��fDL�D�(�H;����|�)�(uZ�5}����U-!z-���\}��k8�ws��ʿr�c*G+Ąioā#j��(�Y�
�
�J@�z"U��/\A�_8���̻NJ�U��]�~[�)"�<�Q����s�㨋1�;}	ےxT�SRF#�mD���^�����^���(�Q�����iF�a6����c�n	_[q]���ƃ������lL"c������T�,6�VM�n�Rx�;�%ph�(ڦ��o-��y)ո���^���5�X�i���ǑğĬ�EIu2K�/���N�b�����~���Én�6����m�s}a>��b�,�y��2�㮽= �c!�e��vB[���Gg�_\迻�a�v�I���b�L� �5��y�tUeW��	�f4 �T�wB?�ة�	m@��`�g���U�Z� ѳ�χ�d�_^��]�W����ϙ/TԺ���otr�g1�����,i�٩>��)5�`��XҼ��]�!�����93�j,�Y�.��g0�榚�*�/719���}�W�V���[�4����{�	]���J�UF@؊b�%dy�k�����F7�k7�B��/�m�e��F;3�ep����= U�bm�4�R,��� �x�<��!�9� عǖ$n���Q��M\$��é<4\��T݆/r�S��:�����@�qI5с�����w��}�L`�\�U.�(�h7���Cn�ϓ'�/g;�(��ԙr+�i�(ʵ�~�G'	iх0�����[ {Ҁst{w����m��g"������ѫ��Uc��u���F��[%!S�fh����g��Tzu^vi�/{�P��mM$���W��o<���(n�Tz��d�1�2u��[�J�:�#u��8�4�%����9K�8zU
c��ċbr'�b�W��s`���G2G��
,e�ѳVד�R%G$ML3_D���z�G�#G�+������:R5"�*�X���w1\�G$t=������P���@��&=E1y�[G