��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_�}ܛ��.��i�F~�~{�J��C�a��K-?�<�>y���yewY�&�_��wr��� jK���w��C�Hxj� ۞�
P�D
��6⼞-E!F�|�'Q7箎h��߭���B�a񻜇���<$��޳PY]�[� $���	���5|`��G�o�Κ:>T�W4��<�y��!YtŶ�/�>W����`y�̃���Bp�2*a�4{�Mg�0�v^n	��b�XȌX�����H��M��TW���ރc4�{jW�-���j�ëMc�zf���w|�*���"������3g��4Gp`���K"�s9׾������M"G�iC(��_+���o=�W<?����y��m��Y���/nv����6�/'���|��wΘ:���,XB�{���������4�Y� ��x� Cb9Z�	P]HY��W:��[�/�2g�n�L�AT��B�`�@�O��U3o��?e0h�r�!9db�b�G繠�ׁ-X$A�,�E����zQ8����L�c�uX�� �;a}%m�`��l�����,+
N��a�2�WY�Fqj�������W�9�C�%���#V�.��P��C���٘����9't�Y򡺃Kc��?�F�Њ���q��6� �� 6��/���9�a�`�lә�<�P�ҋR�ӳG�cj=����@����Yƨ�=e����38\�Ȣ�$`��be;����j��*�~���wQ�:��~�<r��φi�]H׻����^( �ܨ�yԭ��c��[���KXӛ����\X����in˃3$�s���lG��::�/(0Kt�=$��% ��%/��g�)�^�O���I��骄d��m=UI�,�<)�Z�R#jΓWfi H�cy/�0j����j7�#C��>b �eڄQ��OÖp���y�Id#p���a���ےL���D�buBr�W�A�xճ����l��4}�h����|!�G�~��E�jI7c�eJ�+f����2'C��.O���bCc��J����dS/9�z1�b�.v5ka�ή�O73D�>�2Hl��Sܢ�j��:���!Qz�3�֗�L�Y#�K���I=H(kC��>�����e��3��XS�J�V'[�|�������m[�v�����Y'���E �0D�IQ�����rfU��>�'�B�d����=�l������츁$��'�)D�S<=3c�@��Ý�9ua�2��B�埓^��3�$���Rg��V)�n����l�Nf�{�**�q��V(��R\!}�O�tm$�k��4�'8ߖ�p\L�b>c:��߱��c.�Ju�h��x�ye˅�%�J�vKJDX�3M��1���%��n܅7������dw"N"�������I!�Z-':�3�X@����Wt�'�r������R�qf%X�i0���U����I��Mq���>m~���K�	�8��8������:#f��ܛ�u�+�qjWQȗ�.sX����	vT�|T��!͋GVw������%�v�p�������1s	�9��]�z,˝�m�����	#&7����+	/L
�bu$�5b��;�5S�.�{-K���U���Q2G�Q<F��ۆ���v��=F��R��N3:v�XnkŇ��ܽ�Q���j�M��������V�V���<�Dh:�h�i3�J�vIdJ��z���Mq&��`p1R�fn�ť��%%h�Sgg1V OՎ�e�]�aX%�H�?+�|Z& ^��U�Ϻ:%S=�j]��w�D�Șũmm�o�f@L�Q��ּ�Χ1�XK�T��i����@���&"|���.�)�[�H��!��š����!��"��Fd�T�����%i{�@�9X�v-C����ǻ�|~�B1 ((i
�V%��"��9p�tA϶>�CJ߮�>}�&�i}"���֌��u�~d#�!	t�������u�����~�h�N�X�X��%�������wiJ�	��V-�m~�Hj�[U{��p�����UUI�[����?C��..OT{���R��܂�ưG�Ո�_?2nwM*�+�.xX�a�*q�X�,�	��_u"�a�E4PƜ�4�k�/���!vh�� �zC���2l��P��S2vc�w��-��	�6�\��#�IY��U��1I��p��CZ�ň�W��f�7@[l暖|s��)�/��:�*^�\-#����x�"\~�S�45t�1q��-(����y]���lFI�j���-e(I��5x���q�Z�(�`G���A�,���5���/�{���������LJ����ӘӋi��kف�OC�T>Im�J�߀@ף p6��%�}�r���-c�Q�][U�T�gh:K��d�D>���:+�����w���xɠ�0�`E�3�k�%2mЖ�Uw�ku���tD����E�%]�^Ԅ�%�O�7�fj��P#N��{�4ө[�o�<�9�E�3��<�ƶ�G�s_�^;��h�H��Hd�3����\�՘��C�FޟlO�2|���r�b��fi��'|����F�%S��j���Js��`p����r�&�X�u`��ee�pIp��c�L$J��r�� �g�ZE��~e/�cߡ�q?�HTR�n=�%�V��MTb@Vm�;e]�}Z*��*�?�d���Z~�0�X�PNth��KI�Hk1�Q_QX���t���b�ƃ�%]������1WCC^��Zg,K�?�'��t"���y��k<��
k;�����ҹv��T"��?���K+om["�G�ׯ��N�9K6w���h��FC�� ���\dX�XY�ɔ��8<J'�^���~3�ɴ�n�������2�i ��{�Z���.�$�)D�5G��#��i0�E���@�o��S�G/?�� ����"{�(�ρ��>b�m�	cۤ����[�H+�N����O��G֏�H�y����Q[�}��̨[by&8GHta8`�S�OS5�	b����8�;r��ݺ����e,�15��+4AVJ�^�B����fH��Z�o�M�IPoC88������9x�zi@�"��{*�f���7��<�^2P)��s�s����b�}��*0?�v��_��4��r�yJL�Z�����e�&@X��������B:��O�p��+��z��~<7`�J���xyL�ٗ���$*�s��~ �R�/�'"O�������!�Ҧ�0IC����O�T�bA�Ni���/A��c1�cp*&�dԶm�Bz��c�0=�F�;����܅[��ɳ~�J��.��"
�:����H�5`�#*�|H��jm٪���)�N�`�>6�Z��9��[��w�i�Y��_?2���}h�܍\�k.��x����V����7Q^C��*�0�>>uF����lO���3,?���	�����fZ+��(��)DO���5��";���[�x��X}��|�yS��S�s��	Q�p����B��̏K�<����+:����Q��smy_��	��n�d4����B�n�L���D�e�'�K�p�X(_���A#1
�|b���^��i���&ᖢ���PȚ
��Y^�b%W��B��E��'t^�>�*O�m��b�4�r/�����Ufn���J���Q�4� ��V�g��+�_t�|� >���"z@����P^eЛ[�H��� ��U� )n���@!����+���Y�~�Q0��E�8m��ctSi���{c$i�w�Ѭ$C1���QEF'��]��nb�B����.��ߦ�86�6��c�ޅL��$6ހoj��{�]F}3OD�'#T"ז-X	%X���x}K�p�kh��ߔ*v!���z�ى�J��^덋ɖ�;��% �!KIP$�je%�a�z����P���ߓy�Ti�!8�Etk��+
�N�
u���U@��8ʒ韟:����n�r��/,�˅;"TY��V���X���R�L�l��a3|B�B�*?���:��&.���#Z�ZT�-Αv�E9���X�D�	���! ��ϑ��������S��P1;H>�A�}�U>�:����!+J��Q8�M`URd�ƵO��/�wț��8�n{�[u�� �+w	�Mf�Cib懎�4��+m�6>7
��^Qtߵ^�,��iT_���Đ�&� ���[{cs"��ʉ�zx���C�ǀ�ڣ���v�`7{:`d���?�Oa�F����6���h�z���-����)j]���
�)���_~��(#bZ���j���t�#��)_ד��s

S�>�b�W͚
���nj/�E�e��U���0�۵�%��izn����}�ul;Y�ȄB��h�֚1>�-�X��E�����'Y3	�j�E�ITWf����,.�ٷ��J��t�/fB Z;�""�8�����\� ��0��*�25�����\hq�3F��[�"^�V��W�"�D3��"8��\�4]]��i3,R[�V[}��km�	�T���A���0�ig�ļ)PP�<��"�}	�8>���Sy��]i�'�������"A1,GQ���Џ�&�>��ͱ�!�u��~��ASW7������^U�]ڃI��K� <�}�Rk�l�G� @������Օ�G��H|j��2h^��� ��V����х���Q"
ˡwG�~O+/ڸ�0Q���o�P@8�X�B��l6��˓Wz�$'Y������#��q�E�p�ū�Nl}��+���T`��.�7��/O�c�xh�L��r�����{�n	!���H4M��:{�z��]�p K���" �Ft�F|Q��yu�����h[�&�Y���-�s�t����:�I��@�ϗ��	��U�	jY�;�xG>}�\�@�~mr�f͘�$��`yt���{�
���?�S�45ʺ����y���{L'š�(�=�2ּuӁ&hR�,){�V�W.�	Uf���5����SI���2�{g���V��½�~�j J�n|1�W�u�F�^x��:�0rR��!dΥ����Pq�Z�5�(��sI�#�'B?�	����íq�s]�ϫX�O :vb�� =&X�����ƈ�~0����v�b��K�v$|6��+��\�s,�i�@��8ahVw��-[��n0�ܶ`O|h�A'G���[���<vH"q#:M�'EHH�_�s�������𕦔�*<����fd�����i>T������bN�Z�J���[�'d��d"��~b�"��'� ~����}i�^�o�:A�W�L�t�&�Mh%N��@�?T�>Vk�h�1{8g��,����\%��IL"/Y�T�a+j*�+���P5�ܡ���[l���9�����Ic�8�K/e�ON��Zi{�'�r
؄Ѩ�)q>Z����8��|��<<1��Kؔp3gD���*��YKA�36I��4����-�PIS����D]�ׁ#=�r��ї���D��(��2@�B�t�L��h���3A'Z�;"K���D���@��VV��T�}H��ah�& �R3�z}���v��jG�Ab�+x�j����^t�]��$��\4��LV?1�WO�Ӕ����l#m(���~.!d�0;��Ҹ$���?�i��~W�9��$H�p�W��1�'UX�h��NM��/��p�P������Ë�c?EZn�Dᓌpg�T	PD�k"u`z��d���b5�f�-�0�{䬍�.�^kT�}�/6;���Q�Z)`ߢ_az�9х�]�s����3���_�L���ԭ��3�fZ�1��ټ�;ٺ��m��^J�o-�挱i��|j0�Lh���_iw�ˡH���,`�D��4��h����� ��� ��8���t��G����߀C�\�tY��|��y^J�8�_�g��1H�Z����[=����|3��zb	$6�
�;1���-]�̛uF�%��o^�'�5��7�~�b$�(| #�dΊŌm�B�|��x�^�	��Dp�ߞJ=]�\��7���ț��߇W���R�ٹ �»d85"-]g�0�*�&�+Q+P�?���ȡ`�#�������ƴ��{�8���$�p)�d���7v�"x|�;1v���+sF��dE<M9���n�Yj൘1�r'ڽ��zC&��\�Y6J���p��"�`q�^�%Z���ut��E�&[E��5�5�\ �G��/%;�I��9����*҅(�4�Eæ��t�<IZ��8�o49e��ce��4v*�b��5	��ΰ�''W��u>�eE;���$b�T��z������{��pn1������XL�4�l]`���l�vf��M5�w9{	x�����G�|h5~࠲A�D�4�K���/��r	�BrnM�T\�׮����OI�H8�7����)�	���������P��>u�eʊ�K��-,s"Gw
3�2����tZ�q��g᭓�Ǘ��xka�FDz�G8�] ��7�0�Fj�� rOw�Y{��&�cS���m!vY5�qX
�[�P�dL�ʌg�m㠘������v7H�L=Q�i�{y���@`Z�����ɛ�����D����@yB�Az����Y��R�(��P-��ψlbi���#�}�7{�1�u��vJ�ǔ6��D�_-�Fq���	��Yc�i_�쟥����:��++Q�)5����i�Gl ��#�)L�'pG$�O��tQ�G��rؽ6�ޖ�_`K7@sK�wԈ���a:C	�D�0�^���On]�/t����-5y�`daχ���b�H���En�r��w�(PA�*��9`���L�� g�)�H�����U���9�%3��W�]�@��aoF]�rq�:ֲ���m��d��f���d�X�YR����kJa��y3��J�#�C����=�E)�٥<�ױd�5y�d4M(f�q$Vc5��?u�Jh�Xm�!�{~���D���x����lĔw��VnhWRky�bj��H�S\��H�ݮ��(
v��+�>�:;���
O�[nO�3:Ͷ���O��ս���f����Q��JGb�"[�a8A��?���a~��}�;�p��T���@ҶD� ���!oOw�>pu��Bu^��Ӏ���6��#��P�j8\�E�.��ݗ,�����k\�r�וF"]���Mz� A�b]���:��Vt%[�T�M��D&�٤�-G�|�G�q h���l�1���D��܁b2�]���Kij�6�qld����*�
����1��'����K"�Y,AU���!��l��0�@��ؚm���9׏��O�pl�+����"�Ly���$�3Ʒ��Y(��0ΫI��UEz�N��Pd<䈿B��1�C7_������ľ� �i�8��SYchFV=�o����"�Z�a597Wx�l�J�m:qz\��q��ɖR�W"%L�.�s� �5)m��9�s'�a_$��7�iqp4�|K 61�E��@��;A����T�R��TE��� �%#�P��7-�!`58ad�����!9O��\�$_���]�y���1]��B�F.��g\@���}��� �SC*�bR�p'��ˇ�;�E��~���D�镤w6��~����j:=p��}a�L/	��b��~���}��7�=�U�2�+y�ڔt�:g���lt:��6��}�O�I��<͐e����e�����x��ovD�E����� lSЦ�5~w�K_
�|T��~���q�c�N1$�q���l�+�j/C�b�<4'�c��������r�c��gh[Y>X�Kle��5I��Y�u�U�X�������-2��%�ݜ�xcJ�����ӡw;�Ua!�T'����J1�լ�����o�����2M�4a�,�/.���$���0k�wc�&�f�~�gp<Z�w�Va�E�0�>4t���T�:�㧁5`�Hؼ?BZ���LaӖS44��`�[�i,L���9o�ֻ`� Jb���X���m�k�ఁk���#�|ؠ��������(߲`<��]
��B]� G��/�g����V�Z��2�0��K�/~jQ�L���a�Y2��U�c����cȞd��6�G4NP�N�rWc�Q�,#h���KP\��O�> �߶.·]�l�T���e〦*�����L���y�П��`ODΥċ���Gl#�1.�{�f�_��,oiYqMJ���ݤ1=���2�%�#��S�P�Y�gT����7K���j?�ҥ���J~!��ȓ�g-_|l����ȱ?������.�
��(��?'��%9ޕl%��u[�� B���Ib����Ѳn����^ɞ8ĶG������;�=�~@<�� [`Fa�k�j��d��.��N�����!�,��:8�8/����%��6�`;�g#N��oE�����UT��!�K��2@�ZmLQ��FGnd|�F�:�����H'�<�,`% 4_9�	3�����7���Sk��M�����$���Ԙ�a���)b�~�\6O�6%/�(8oqog �G����cbG��\զ�Q���(�Нյ�� �`���|���0���&Q��p-�;�z��,�7�b!�zN�tRu��%r꣪}�C����MX���mߵ�~�)�xr��C� �
�Q��+�e�找7�}��Z�+ή���L�a��D.{���cVrE�2�KQ���Pj�+D>�K!˽Ѐ>m�j$�)�F�@���{��^N����D�7�OR@���0Z)�t9��a%H�p���\��%��B��9Ԣ��$��o��үL���0��;�Wq�7������j��4�?�i��ӝ��&�o9���
K@W3H&�E�י�%%�w+�7��P*H�N|�Ɣ�]t7v����7,���9菞��M�Ϝ�䙑�����В�'�q���� eP	��d�_z�� �R� 8�F��p�Oy%�!V�*�&\j��\���Hf�q���?��C&OAd�:�/��\�ڄ��0��qwBn��1]��sY��lf˼����m���\�,1�>�c��Yi׽���}��Y���{��*�,O��r�qE�Kkd���"7q�-E&������F0[��Y:EB�_\U�8m���X�I��z=�n='�|������U^Ê���>l�G���L_"���ƫ����T����Y�:.��IO�����剢/*�V��&��\$��FPZJ{t�G��{Pӏ�� J˶d�z����Yhf�4rxC�0�3�-5���.	�k�Q�b�y����=`�š�Q��M��]�ޯ[�������4���f�֕�EH_�XV�f���{���RH�c������z4�����Zʥ��]úT�ZD���rm�[�+�f1�G:e6>�a�IS��79����{��b���FY��`�&=���ص���G�p隱��q3�C �xZ7�Z�c�\� m蠵���f��o,5gFl�W�R�ڕ����e��o��x�ߣ9,q�_*�1&x���i/ʁ��g��n)c�4Y��/,���V��Mv�<മ�������@�$|��
Ūa��M��7�n	��-ߚ4|f�<-�-��f[�(���H݉��x��i�kó�F&0r�ҙ�  w�ZKɇn�ZX��h`�jz�R��Μ�7و_��TV��:��5�P�_u���!�4Ghj�15��֚���Ҏ���(ن��4����y�j�1�&+,i��@�qrR��-O�������z�6�b�2�S��%�$��6�.�A��1��Gb���^J�x����t���.aXW���יH�o��ò��z ��Wj<�3���+_5r$��l(s	��̭��ߚ㕊��_��s���񉒢��NDQ���51��-���>�o*#0�%u�DI	�,��1,�~xa�~�f�آu�f�N�4Eģv��2��S�&n�b���,u�԰�1�@b�yw�ꖲ��I��w���x
H�B�^'垼� C���u+bEh���4F;�Ï��g(��A����"�t��3i�9� $���g��34�yc�nIJ֡����f'���
{g�2cK���wm@�eUa��-��1n��Ռ�!C�!I?:[\ߡ�H�8�4����mu���ݻ}���@��J�E$:����#u;��%�Õ�w@-�έx%n�����cd��� �}�b؞�[բ�B{��P�ׯC������O��c˱�՘(�Trrf���y۽1]ٝ%J�j?�
���
!����"a����� �y�����zfzJ�Y7s���iQ[��H!�2 *��k[�Ik[��å�����(ť��`�)2"%M��ŀg�q:I���ɷ@��^R��
d�'�b��Hb>����Z�K_Mc,���C�%����9��|uZ����NF}�d�JC��E߶wi�Rde5C�?uA�*�h
0���5WY��k�4;��Osos,,���ZN����G!J���ӵV��r��A��S�k6�aT��M	o�G�01��T�����~�ŝ����u��ެ��m�`��Z/�_8�H�{������r*$��m>E�k&�t�!uN���o#�:�i=Ofhςb�4
g�cN!2�,g;�/�~t��"��ҭ��
0���nA��u>޺���^Wf�ʣ���c���F�r�.�)�?S��O����mj>��2&�|����s&���g��/6�r��9%��/�$iP����ZQ�!�5�����((�͘o�^���btS�g��+�p��<�����l�w�:n��Wl�v����)��6z��]�5Ş��bB�S�Ɔ�;TK6(&a���>�`ޞL�ܽ	��[l�}�&���+�2jr�5���O�-�'P??�Iw�8X�
��{Gx��ź��(;�&���)bޫ)I����p�b$+�L�J|J�=44q����=ah�c�����$$�H���5n'#g H8�L�����Ldtf%�t����fQǀ�n��%���*�P�� 8 qh�&��K�2����m��~)��y�ߌ]V�H?���^�G��U_TL
�#���� ͒}	;K��H7��;eP��;����J���d^X &�ۏ���̪��W���Q[+2Eкڗ{�;�Qq���KS�(�˔����L.��8���U	L�Q��ej{%��~ְz���-~�J��K3�aE�R�M鸗�a��Λ0i	��ͭ�2�0Ε�!7�\�+���~F:�݅0]�4k{; fT���Z��Κ���8� ��P7h	�R�4f]2믫_��)p}���߭-�u� Tj⠎����V�4)�S�e�R��J�֜G*ݲ��_�*۳����LL�$��8�v����'P=�Dƞgq��HY>��a���08_	�Z��3G���C��Aէ�|��uq�8ث!��K����X�z߄�A��mrvgHܲ����eNJl�:m�#8t�c����r|*yO*�PV,ՇO��L�lQ�4?��Ʋ��ճţ�Y*8*
�U�_L}��f3�����t��;������,YՆ��7��Yu�2xd4TD�����m? ���MD�.���Y��b�6=��}�|�vc�?T��P�+J.�y�aF�ZnGcl�[3"�m�M�@���d	J)HY�1������
v�'Q�gE�8rq��8�w�����oh��W��7��u��)Qx2��t��`?����#� �T��X�#8
���}���W<oAd�h�jo\Y�ҹ�Sc+dߣ#Zw����x�^��#�F�}�d mÚ��r u���j�џY���LY�����G�6��/��(�d�V%=��������	%�v�&�.~ G��HN}Eϯ�����/��ۺ��O�@����㭇�X"$��P�a�2��sgoPS��hm��v�,�!Nt��өr߰¦X��s+_����݁+�Wgѩ�����f}r&y��C��jF�ϰ �3Ͳ�Q�J :������Gs,|�w�U�Lʰ��N���l��$�%����/mP�J}���fCq�x������ ;���c���sp�ٳ��!��K�����{G3�#++�cp�b��W���o/{�QK�/IQ<�ofW$ș�P|\���ϼ��nLu��7��k��� I0�a/�uy;-q{Hdt�?�SM�>��TZFh}d�n@��1m������^Ր:s%5��Y���x�A��yn]��B��|�C�+˭��f�W�� �}k>��������c_Ya/�V*k�j�#�����U� s�\�Φ��$��g��u�D,���v�KVO>	�Ϡ�9��+�D( �����Q��bB����������`D����0M0*�ʑ��-�  ޗ���7J��.��mΚ {���K�t7�s��#Z�	k�:xd�`uQ�0�l2P'J�.�Y*σ�\��_o�ʎ+�u_�i\�sń�c��)�B;������EbÌR
Mh�p��cI��<�>�8{�Y
n�-U�0��.T�q��8! ��ě�+���.V��>���h�U�����,GҦQ9�7%��1�ѹ��`�����.E��y99Ո�N�K����m�^�]�e�VB0`�F��ѕ/>^V[�� m���%�Fg�T�qb7���cc�"�-��Y\i�Gde�*b�P�(�@h�윚��*��E�^Wg��=Q��5�Z���}W����)�v�?�>ͫR�$�Z�Jh}H�)���0U �\�N2����A���tZ�,�oaN��+rH��	��K��0�����];V�K��?w��Z��%��BCD�!�n��BX��J>�a�~�eg�U`ȵCG�Gg]�^�No)g���0~�c�1Q�O��_�i3������+"�2��PlH :�) ��;O�Y��'��젛���6,$�lO��V^s�y�$d+���L�=�$O?�<�`��w�9ƙ�_�M��P8�ߚ�&8�ɢ@-n�pE��Q�2�2q���2����	wМ�t/ �A�m�T3���$]���!��Q.G�>�}۹i��2���}nS�����0���Iw�������NR�%?+�T��p�\o���[7E���`n��L(R"&m�����)�$�(�.5�q=�J�Ѽ�+�\��u/���xM�4����3 N�7�랩�h����E�C*����6�~��a����:�*sΞbq�����ÿ�d�:~�ޘӚ�U��cν4y����D�i��T���jI��)��'�m����i�����F�����>r�ME�{��\P�Bϸn�i :	��*�N�]���n� �p(�c�*�	*P�"��l-���B�t=���[�tXr<6�.=����d�<QIт��hM
.M�Z�h�c	����4�П#dOk͐���#I�P�PI��2z�R]\H�]v�<; ��O���~���Eo�yS�,�R�-P�xv)�g�	�7C�¼�f3'�d�զ�A�~�sS�>�j
LN|Vi����w(�F�Q[7���j�WͿ��_�}�8�G�ueUSD�/��֘�d��%A�e �P�IC���<"��~ơ^d}&lF����!?E��3d��Tr���p�6��gn��C�t�6�B\�=nw�d�f��QJ�'rP�`
H�����v]ݓ��m[��櫣lف���$)�~$(,�e<��`N��%*�Kđ%�_}�>
� ̳cf�3�V��\�5ݟ�"6�P,�	��8W��L���Te�X��c6��e�o��G��5�P��o������(�a���-�؄3�=��/s��e�U����3��j�IS�Ic��{~#��{ŞV����u8���j�cN��%�����*��jVF��Ό�T5B�����Jc��֮����8�ϹEh�G��]�&(/����|ΰ'om�u�tQ��͒cP�sw��"�%� ƎC�wC�f���+} ަ|����w�!�����\��\��"�32���.*N�%����M'�����{�c7��4���ͣ/�7N����H��������5��tq�r6]ы���cJ�/�N+�N.lv䶄+/L���c�ݰb���]C0.S|G�ר��e��QQ�m��;(A�.�'�x�CČ,��j�xF���˸����
¯��������.��Y�z��w٨�|�"�%6���g�=հ������egx���q��9�B�A����U��:����w��
��-.�e���yT�����2�
d���!��h��� d�S��_�W�`U"'�\ ;�{�[�?�!벉�u���gL��*��!'�-}:�+:��s