��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ���\::��@T�qRk	v�z�U�����W�Kۘr�YLZ�[��Zwuy��oV$�#8�N/D\�ڤga5�^�F���,s��#��7�PU#����a�$8p8*� *"�[[�C�����O�Cߘ�m.]��w�L}��dz>�~���/�{�v$��|ʆ~�?O�p_�I[���Zc��-l�#�ª��dwz�x����_�7  Pa5�5/+�U�<d,t�H��Aҩ;��ޮƏ����p�����K�����4�źXWWP������T+#i6*��ǹ �n� ��'x�c����y4�M���ʗ�αt��v�TT�LD�X�#nCM>	v�dM�}��X��R�>�Ǭϲe9}��GҦ�f�0�j~A�cJ8|�2�U��\��Af�&�wM�k����'����p@5����'������ɾ�α���G��\����Zo�1���B�Y�g���$������n\ ��4�[U���߭t�eܯ�l�]�k�hn��[�"M��'	�x;[���"��b��=YF�8@m桾�vE� �S.�U�)�d	(��'�JK��\��q����S������0��&�pP�\d&k����X���4��@��]���E����Au�N�W��^�\�U6o�'wjb��2OS������L�z%ET�Z�S`��tK��1�24��As�\��,n��柑c����=��0B<۔w VD����K��u��)T�\[� Qe����=ڱ�-��,B��R�>Od@��7��ȳ�^2�+=݈��4��h�l]
���?:�	*a.#*b�����r�5[�$���eIV�k�����kXP��3������ǚ B����B.e�m҇�rџ�϶�	��I�zŸ���&�F*��M^���C��	麪��;R��-KM����څ�M�/�ͪ9�ҏ*���S���Ǣ���x��n�m�3,T(����H��P��ZO����?\.����I){$���G��i���*����SuOOSc��	�ߥ����TNgz��l�x���ʡ�����?�}8�M�|�Y�����'�<�΋��.�vt�|�>��֚��"�w���w�:�w��7�M�nC����S�����V;�����;ټ�]�J6$t������wD����-���S���7��ʿ�s�g�4����[����oˇ���e�$ˋ�Ʃ�ݓ�p�D4����B��`zk��� ��93�mg5�Y\����4l;�>�����a��|'$ݒ[�M%�H��狺�}OWn����1�U��_�c�j�������K$���Q����u��X�˥m� ��6�ʪ�*~��j>m@�U�����;����O�J=8:�@r�I�@7��u�]D�((�5+U��6�=��+� ���h�/�_����=l�:~+3wj�|�]�2���H5'��L��֖�}�$��]#��#�{<�+�s`9*N+� ]�aCÒe�/^m��`�'G[L`�3�1kV-�)�U�8�υD��!L�Ms�����B $�!�x��+K#��ʈ:1Uė��{���WJ\����Ɍ��4��wV������
�}� '?f^sȶ�*O��7��zB��1,�X�2��A�n��{Z:B)��A>0�Q^���Bx5���ސ��%�E����Ҭ�s����^k���	���|o���"�էa�Y|C7q���o��s�2s��E�a��T�S�>��ґSAv�Ɇ�[b"H�.�$��;�oP��EDM.m+ O��T���=܎(r���e�̟6]c�	�r�z�73[X�]�}���?�D_EHi�'��*T�z��J%���W���r�N݅OvR=L�
�43T���Qe7��\iҁl|���1���5��"*,"G���BK�%��Xur.���v
�q�~C�k�)��ш�24��RB�|��A_���Y#q���!�\pp�se�0Hظw��q��|�tL�Z�PW�n'�@S��޸�#���d�H%Fj1J��kE�Le H���2��ů���#.'�=m���!�
|���ӧk���d��vί� ��8���j��wA�:?�(YLC�{��UiS��G���t��A"<�`Oqw$�����B4���+x�FC�Sg�8l�:#�s��U��_Q�ſ� ��3˹P7��M%;�*��D�>�8�"��d�Dn�r�?�*�j���5k��'��>�W��z.��2�Y���(_T����0�4�}J��[�a:���f���ͤ��ax<y�Yd��5_�;�"�!�;�XN�<�L�7fcJ�e/$�#�6�3���)x�F�tĈ�
#H_̼�G/��WI�i�*�_ww%����"%z8�3��ǧ�p�����&�U%�-�̘0�g�o�3��;TL�Hwz��1�X�� U#o����rY����~�ޱ��xs�U��J�T��N>�����ϗ�����2N8���C?����a��m��X����(���׮����	�g�\��ʲ覾�}O}���c���⡐r���?KO�=G�@���ht�{�d���U)K�h��&��|YY`�|�#qں�[����3�2����(ޢ�vZ��5�B`p��=�u�()��h�hz.�A�c�kcX�����fwQFW�$/��i���!�&�p��6L|T�u��Z�K���7��gL;�4�Ѳ���CT�2���l��`[�d�զ�8�e_G����\Χ��f�rS��|�IlG�����4\����, �׵]a���̠%����/����!<{�� o���;C]��V�8E��F�:⠊^*���!>�,�'�b�k����B�0��ʍ\��?�0�֚�};�x3��R�뷲M0K/(�'�e��4�D��h)��m��4t�K��v�o#"Q�i�4�8E�� QJ�򱩺r,f�e_��,ĨZ�L)mĂ����륣���#��ݼ�Q=�����wf��T�e,t�L��3�tS���Kkg3fZ��C���c#Z?�$�;��w����:I���)����� �]i���I��M�[p#F҂5��܀D]57�i�Á� �T�ۅV�pK���^�-�eqw��UV�缔z�(=>���,k_�.�ev�-�pq1S���)�ו��]��T��W��{��}�`��b/6�-��)@Q}΋���6��*�n��3�r2��*�?K)Lg�H�$G�)E���7v~���Vʉ�E��z��m�� �0�F&�I��"Z�L����i���Ȏ�\$���&�� #�sƧ�S9�eV���-��t���O+�Ψ��#��?P�0���[���>�NQ��5hܙ��Mg���%�w�z�9��^���/>3�|q�@D�/� �2�������3g�j;��݄����$���ي�(��ܥ3��CS�HGm�[ ��_lT��Ȫ@���-��/ӏ��O
��e�����Ar4�5����(����^b<��!��GJ�|k\!�|�&�>h������������tC�f$�{�_�u�(%�x�h\�M>�:ai�#m�c��Y�g�ږ�z�f�<C��+�2���|��z���j���d�i�:tv|������r����z�B�$c��
��'ێP)�MB�������^�q��PwW1�P{Jb=�GZ�a"/��0�x�ɢ���t@��5,��n��L*�x����m�(�3�ry���h]v�۶V򉹯�g�z���` ��#��~�D������$$�N1Y՗��A+5W�= e�>��l��5w��s�U�/5���I����� �;��uI�v1�h�4'F��X�
���,�u�/wZZ&1b�����D�l�	Ռ��|�b�v^ ��L�����&7��.�A����(ǆ��>c=�"��skΛZ`�#�F%R��x���<f@�o��S�pyW�0��N<r}�歔i;�xᯜ��i�'�~<u�c�C��-<���6��F��o���@�c@�	�_<�����5�ܙ��?�2���NLM�x�65�Z�Fzi��d�o9�cМh�u���כ��L|�f�Nw2hؗ���xכv��B�&�)��b�*�"(��4�h�:���F`~�������Qc��J�~�\n�t��ֱR��{Nz�4b���iVgÁ�F�ˆ��O��Z�D֪�����
t���8��g�͎1';�1�c�Ϻ�.Y��.�"U%y�~+�����[��xT��>+�l�1�a��uEW	�6;>�:'}��{�607dpHt�t�삣z�^_�(�S�,�p�xY��IW$��c��k��Я^�������n[ ���k���B�x�E�!q���F<T���z?Z;U�9����<x�`!Zw��"�?�"� [V�#��|��������pø�n]�}����ꇖ��l@Q�}�[�e;"�c���[�8Vh���D����u����8T�.m*�����˫x�� ��@W���!v) G�GU;,%v�G��i�i;W����ca�8�}������[�M8�wY%�X�C�5����=#�{9���o���dL��3����E|RГ����X18�_��jWC@�x���4ޫ�������c��؏erV?0� � p����s��@�z���d�o�'�`'�&����K�Ri���9��R'�ܐ�V~8]�l�˥lE��Ү�0���;���'Eu\%<V�ו 9�k�}G{eG��9�X&��/]{����Iwy*��
�e��fN���v�z���Xqt#���ɢ�D������/jw��pp�5�9
���b�u���ú��;��p��#��LD�3�h�\� s�̭6�[���Q�DB\�|kMF��Q"�X���)�J�O��Zr0r`4y Q�"���N���ޛ�R�`L�Ow�g��Z-JrJ/�?�V��t��v�\}T�pqV�;��q�.��G��q�7�;�Pc>Z�!�D��T��Aс��rY���8yE�U5A^l#R�	Ϩ��3?������L�췼q[��������C���h{��'���y�Q�[��k����#�ԕu<�$�ⲻ\�ܖ=>���^�&6j����:)�.�*��Q$���������c6���������|n��������G�/&Yu�N[T�hd�;��lI��ޣ�Z��
7WkȮ2}
 �������:�\���<	~�M<���bT=�$֞qE�[]����Y {���K䟈F����#� R��~�5����* I��qu�� W��H�kQg$���,'���]�O��^I(�(Ȯ �&���!a�5:���1b��"����R�ewOV5h� <7:}���q�Lcj��O�,��ln��H&;��}���e��&ǰC ��/����ԙ�ތJ�˘�~}��X���#L�2�)��˗�}$��|u�7��E�98 �\XIeU
�J�R~�J����L�kg�"��'B$#�g�k�H��W��pF��@�<Y������R���.��E��=w�����E3BF�L����dsi��z�^��}<�����U��KĚh�D�%7�y��|(5�u�z������?JG����>�t�nn������Aݰ�]�����~�l�>�n7T�\��	{s$@�����V��e-Frq�^�����I"��e��RG�����D�$��v���b{�sJ����5�V;/n����[���=�=��@�.�~�6\���?�K��s���h�ĳ%4{���p���l��J��+0SMj�{����!��ޕb�1f\��@Г�ͦ���2%�QF������'��6���]55��wj* �Go�"�h��җ�U�<=W���G�S���!^�|?���1�ڡוް)&��%��o� 8� 9�W�jk��/S�ex�Tp�z��6l��8X�+��C��zZ��_�f�8��3k����YR�ԌGT����K�~�Z��w�������O=Q�|��s���o�&U&~4���@�!�wX��e��7/�eu�uc�d%e������b�{�ho*=��Εt�'uz�����4d�ÐZ������}�X3Y3��͎"��RH�- e$e1*�G�����r�� b@�Ds�e8v����7~֍U�Lh9�'�.p~gnt��^��RP�}�mč�R�r��u@G���%����3�L�\�;}lJ?����R�ت��͛�#��kR����(7�'&�_�@�M��6���-�s����l%7gh�'u.�ʦ��|�z���29'��p��O�h��/ "��/]
�g�����ېd�g�;\��0s�5P����pַ����og��i��V�FAcխ"v&�N���$. ��Wy�D$u%+�S�<���K�3p<\���M���*�V�Ed��[��$��I�j}���qBD��
�pPH/��\�������4�����0���Ic������󬲉'�A��Kzu���0� �`͏���R[+w��2��5���r��7�Bp�߾�BT��+Dz�W7E47�7������~,(�L��OZ�ul�Q/�0i�@�q��Kݥʳ�%Y'?��̫o����@}\B�����YW��N���_�:�>#�])���~����h�~���>{�q�Q��j���E+�����6��6GO��)��7���{	̦E<���m�K2��1�Pl �II9�k�ô�q�(�?�x�Y����/����Q=�mh�L���|t�zޛ��HE�|�:٤D�V�1�TX]I�q�Q��5���IZ��.�N�m���(1l��@)-�?
�����l�ie��]^�H��E�(|���ZT�9�&���-	�o�I!ث����ڬ�i���F+ |,�繏?�
C�
Z�/��r�~��� �����E}��Ϳ\��a�ke*��s{-,�/����%�>oH�ON����8C���9wN,��^+M�+���F�ޫNU�	G[��&>hR���J�$>��uJU�r�\�'�Z��6������]���j�J����ŀ��	f�nh�����[��ׂ�G�G���,7�Ez��9d��8u0%t��ekЍ��m�#b<�N�`*tfh}N�c�TDwy�c��<|o$�7��
]@�o��2�<r�]"]����+P��oG�h%���lH�{d��6��/����w2M ��X�F�z�J�Q���*�tm2��j��ZG��B�GM(��������4-�����ږ\��q���P�t0,Y��<��lƬ�ڕz��UP]�*��?�I�/JwK��f�9��w֋��Q��+����k����!��5\"U86�rb�S@�{� �����2�k�b�Y%T�؄���@r{�l
��ۮ�)�Wǯ���������������g+��ݖh�G�jtM^���n<� 7\0M�����Xr"���k���;q\��[,N-c5��Z%��y�c��{ �!�,��Rmx���c�u�;X��Ѐ�%X~=�V�J��
o^ʑ2�Ƒ�P���ؓ��'V ���L�C����<��Y"�_�Fm��Ŗ+:^��,l�5vvA��S|��7���8�0{��#5�@�Xhj�(i�k?z�eb<���s��~y�K&��J���&�J�>���*���c�\��(��o�`)(1K�a��}���x��b�yf�Lד!P'�y�Г��ǟ�k����ѝv��'�A�S�@Kp��"�D������֍��qb�&p*4L_Ϥ�A���tPz�/�,2��y�h���5/��[Q�_#�/D�"�_k���o0��D�N�N�O�)�O�!y��N��TL�^�]f�Z�Nx=�G�;����0[-.'���,��αO�,�6�v�s5�/��P����9Ւ�|���d�Y�p��W�
����z��`CHBb%,�q�@X4"رw�C�I�+����/Ϊ>Y��-�ia�X���ˊ��������RcHת�e�zb�%�*F�\I����IU�M0t1&��&��V�:��IY��[���Hna���,�ļ �r���Qw�����*NA/ygv��=�#@�b-r;���UrIʙ����[�t݀W8��eع��hm�����i��a�k�����k�(��0��" *@_M�}�zn��$���?B� jZ�[���;n�y�O��'����@s��``� ������*����ǕI2qL3�?zQ�=���>��ذ���|̙�!P���]�y�!8���2l����Ra/�d�KC��)N7y��
�Tzy	$W�Ȃ�	�,h��Z	=j��^Dt��UQsM^M��Ļ{���x�� ��Q�B> J�l�9�	$��m����|�������r�0��X!p?� ;�B	��ҳk�B�l4�䣂�� �����!�[qk%�]�yH�����9�����txx��g���3�щ��p�A�r1Ҙɞ��_�~����I�r��-*q���/�u�ɂ�զÓ�o»�o��[Vb�B-�c�
sGpΙ�H�3p��_,q}qQ����xh
��f�]������/RBT%��0� ~������\͛�|ܳo�
a��X�Ҥ���	�3��(�
��9��T@�TB�*.st�w��.#S�:n�B,��O����&���>���
w$�<˕'�Zlj�������@��,Y&��˄�+�e[ԄS/�4<���*�O�F5]BAJsJDg�cX&�"�+�a��t����&Z`�d�����%X�.����d�0�b-3���2-ё���e#d*��˜������4�s^O�0�!!{.^^����D�@p%����_L����J>�˫|�d�oHS?��V��d��[��:��ܛofj�v����IiH:p)z�u���;ȍ���'|��A ��_hq��S�����F��:����������+�@���L�Fլ�_�D�g�}�my�|�TDY/:!���($�!zw�~��+�����4���\A�rAK��3��tiV�ʨ^Ӓ�ݼ��LDP6L3��F1�oz&F%�d�akO7@��8�G5A��A澾���?T�~������!h�N7��ʟ�E��f���!�l��Z�gl}J��C�XT�j2�&�U���u�����ب�ds;P�᫼�#�A�mc�ߖ�s�����*��ӓF�#d�E)ϱg����AGu�*�p�f �� ���j,k�NJ���.J���i!�]( �Wz�r���j���2�i����s��|��<slw�n�/�Ԭ/*�2�f�ak&[e�n����;no�Qݦ
�ǳ�Y&D}�ƛ�R&��(�fW�	�]I���E����1���E�m�-�b��Z� �~c�8�p0�,(28ԯ��L�d`�z_�(
fxM��=nsCե�E"|Y:�@q�y'��`���H%�`���ѰP�m_Q��r���2q��jܐ�^)��&g`De�g�� v�Er4b�('�֚��a��gNiaϽM������!c�~
1�_O�;`���p��u���>#�����!�����
f���Bzzs���xZ¿�X��z�K�v��*6\>�ß���]�9����0���5�+�7=�XP�j��nL}an� ś�>�a�~���X#ug��{d�{���I=�8k�Y;�l�D�􌙉L�m>�_��U~�^�ڰC��+��>���_��߯�g�ԋ��3��R�d�ҹ�S�V�������JW��z�0���ܵ|f^�F�f$��r˺���_��$@u�R}~R_�T�,��H;����!7c��n�� �҃�úW�x��*�� �>]J�ɴ�g�Rk�Oߟ���U��&����n�]��%�|����`2��WȂ��G|F�%��'%�1�E>g0�:H��W�Be��B�0;���������Sj@'6 察��^mpj��bs#A!l����]�� � ap{e�5b�[Mʫ�{1[�_���43�v9��̒1��Gb�A��\�R�kn� � Po�I ˱Fg$�Zi����j�t8�{d+���dHG$�܇�Ϫm�/4��8����eb��{|on�%$�7U��젣0�Y�(�g��
���2�>�}�P"�k*�&!7WK��˛@��Tk������T�z���x9���X?>�k���(u<�󽀋���%f���<��V�t�[@D�?Z���w���Ja��]�cK����}�P]�N;�~@f>���/!SLE ����Em�w@*�N�H1`M��TK]W>Je�����GM�Up%���R�6�S�H�Ϣ�>�̆����yuj�i7��[�b����k�����B�v��Z8*Oc��`�'��Ң�[��V��YܷdƠc��U�kj<&�I�/��P��h���R��p��l��e��R�a�1���P��2�).F�F�m��59�EI�¸[����#��|�09�#��5�P�Z�^IS�y�x1�iH󦢛�3
ZK�ts�ê����Iq�Q6�<����h��F[q���a�����{���B��S�M��M���3Q=��\�]�u�k���'=���O��$]P�L��}N)��Wҙ����-�e�'��������zӣT<-J�fN�8�S����T�q�������ed�X�������+�r���g�/�2Ȣ~nN$���B�=0[K�6�3��w����k����l�k�Ou�d#�ɟ-���K��D5�:֮D{�O����F�qZ�|�`����*�(y�H�.��0����B��9)��]l���(�FvH�'����-� �,r��"z�J��l3Y��"gi�v�e#�2T׫����v�΄Ğ��`�9dSFfQ׏-��R����4($���� 8ި���J��U}�ӥ��+H����4�V�/�)�
�d%{��+4�(	T�0�� D�$����(TZ��=�H��	c� Í1�<B����hY8{L�����pK�6���͵��=��Φ;�F��L��2�8�?�1�x|sߡe,�ͪ�{�I��O_/w��ծ"�b���+m�7�0wVk���B���y7��0dG�Ժ�b�X�W��P�e�,-hi. �F�gn��W�xN_����E���?���M�KbD��6�+8��s*�� ��L���m� ^n�@��zJk�k,�����Ů�|E�+��� w
Gu��>�?�u�"�']PjlS��}���l�Gpn� }&�g6a���ٻ��߀�{cX=�h9�L��t����
�`�D��ۤ@{<��?�eG�����74a?�o��y�{�+R h�Qnk4�/P����uɎ�w��4=̊�P�"p��4/��E�Fꭱ�T�;���x]ǁ���-;l���ԅ��\�ẁ����AGZ���'v#x�FM�3uow��Ad̮w����Y����#n|f�B��ȵ�HϿ�:*�tP�j
�5@A����B]�*6���;���]����G>!��?��΢�()��θ_c[e3q�H��1�>4��dFV�m���c*�)�JU��JhS0���u��W��@������?�_T|�N��J��&#u�Yc*��UL[b�PiM����5.�3����x�l����rEѹ�c`�v8�i��ǣ�W�(���Q�O��5�F��v����8����/��t���Ǳl�DR~	<|2t� �A�;�<š!�>�^]%Ǚ9�l�`m�朗U?�2��j�R�nX>�ط>*��K�
��R?2{gQy���C��Ƭ:)���+�����+�����	��b�Ч��&��|�oўѿ�Z��H�a�@���o��M��� �Ŷ�y��yTu��Y2=��w�&a�8:�G3�l��#|�Z>@<~IB�u����%\!�~]7q�C4#�pG�p�\��@^u���~�<s�ˏ�Mw�w(;��x�CMG�?N)�UǭF�tWAqG�R}Oxʩ�(�d�C=�����>;Cߏ�&����i;V�$�&�0O6*+������E�q�=X���U~�sR���󇏩ٗ�����aK�f}e���U���	�y��Ϛ��J3�JMż�z�z'kfm=��c��=���s]f98Y�p��˄�k�������Z��a��ո"\���Dw~r2�S:����k���&+_�u�G�t��!�1"�:�i��eF��Z�H��������t��h�@��H�����z���u����M�s��/U�s�����/�~.W&5ǘ�S��(:��M�yrX�1Ŷk�o��s83��A�#��A���2R��5<R�pR�T-���RY}�=���,|��	1|X�O�	h�~6>�{�Y�y���"{ �u�(�����c "����m@��Lk�L��i�,��~n�D�vJ��{棐�K������Ƽ
%��4�m�Հ���˳[񆗄F��`�.Ⱦ�B�����R5_i�;U��HK���m?4���aY�K�[#�!=i��ϣ����{���,�e���{?������}z�/�z�(2%�0���z.�� �O�m �a*�5����n�+�$Ǧ�|DB���!�[�X1#9��8�k"�.׷u�+^�
"m���(��4���6"�H�����f_]�����k�$=�����x�3�~�N
~׎ �5��ѸP^M����3�-oM�h�̱��>�������A�&/O��S�p���k'mW��,<��M�'r����Ku��!a�[Hc/�����fU����$���nڊ�~��Q�]1	���G�K=P¼�9�;k�_{	۪L���h`m����"�
SF����P�_p��
� IyA�
Ic����V��FM���Q�	/�T
�R��D"٦��|���uE�,�
���;�k؂�?����4��/y�D�R���U��b+\쉤{���ҀGV��h�-��� ����7v�[@x+��X���7G�^Bwq(�Ps�D���mCd�_Bg2���O��p�/L��>�z��f��E��dj�J��_3����_`~��x/^��h��KS��Y��m~�Iv��ş >/�r����q q���4Uy��D
�z�0 �p���$��i>4ZR��������oO�-P,��P=�2�*y��G�Q[Y�\�Re
�ݖu����OԈ}�� ��DO�����34;�wC���x��4��-�.���jkڠAר��e��_��uĆ�/y|=^AR��!�>7���}EE��rO�Pc�gHn�sE�U�$0OK;�GǮF:�+��W.Z�
QF�p�Z� c��GX~{��%Z#\���nk���(��o"Rз�,��<�{H�9*����̛��-��cة��&�C%f��竡S5H�������|����18|m�m��ĉ�c�g�����AGn�];O�5���ݣƣ�D=Zqt������3驂K��U��(ys9�M����Չj����ZN�������8��M���7:�j,*�I#[��vy�d0���+�ڃw���/�����d����P2���.���"�o��d,F��7� iS7��v��� #����c�W�ï*I�٭��?Cq2��EsFK⹃1��R����k�D���x��ޗN��=说���0㡂@��@�ҧ&�t\f>��Q)������u�]�}cGL?��[�a�i�iv��s�P#Tz]`�2���e6�&�)o� ���U@g(I�|�;�i0.W���;��Ø��F�����b��Ȅ�E����!E�$���-[݃���d����w!$2�/�0�n8F���b�U�weV8�97n��n�@z�� ���>��-q�����#倒�,�F��n�(_E����X(�u
A��uf[-+_�vlj<B����˹����&>���=s��Ĳ6<JPY��`�f�D����zY�t��L�Eqs��ڄ���3�S�.oZt'�r6A���ǹH�$f97�����DC��b�D"�yv׉��.����S{:�R�9!_�2��ސ��Á�����m�jM���њ�>�S]�;�Z��'� �IL�Z�5@��.Y�J߬��S�@���i�n|�����N�=d�q��S�E���5�Y岷fW��r�j��{����i�(G�އA�� k����}���]���D��s�?<f���nHڷ�Z8x%���Em%�zf$�D��yA�rt�a���nQ!�����cb^?Ƅ��[�)���sG��,]?��:���c���ͦM������rZ�R�.A�����I����B7g�XQ���˳+�i:W[��Hg��:Q$�@fy���. ��+g����mE4Xx��(]��W�3�Z_j�>n�X��ɶo2_�s��N!����Z������@��k[	���cxh�"��(�� P�=O�!0�;�q*Y�e�[J�ޑ�3��cO���jeMFk@�i_�.�<�g)��	��q��2ٺ��(�����4�;�s�]�>�lD�����m�k-���5�K[�{R��s)����V#0�i���b�n�m��&O�7�{�&@P@Szg�h�I1��f���JA�N����±L�zd&�o�"�Dg�����˖�@{�5�(�����F}���%��|u�I��%yT��lW ��iI��'��dl#��eD�炦*���.{���(.����������R��9'<��f�F%,7N�HI���!G�t.O�3�م�"��\O�$?�pD�A �Q-����?��QB8�7�k���<I��C���wH*�J>�`K�2Sgl*�&cr�mC��;��Q�j�@�1m�՟0q���j쪊=����Q���ɝV6�w�(���y�:9Im}�t���Dk�b��4����Ćpk�`6���A>w�x
�� �b+ d2BM!�;{��4���uTLE)�O���G�ݘAm�Šox��4��5s!�@��)]!�-H	嬾��sM�s'��kv�^�g�,�ل�����;�;��(�a��i�a2u���2�λh\y|xG�nV���c��듾�!v��?���Q�=�.�<$}RU�����X�kE��n�k���P��:��m����v�r�t�Bͻ5pB�|��w���+����f�7׏�]#ċ����I
�����D�b��Q�������xѝ�h��6:��L�Q ��
�gC�56��&�l���~�y�'��� �x\й� ]';$qIA�z��j]K�f��#\ߚ���g��y�yWc�7��I�h9�|�:� a���L�/XUҍ!NA3�ulQ8ƾ��{m���$#�r�y�O�j�.����{i�&���7%��W�ٰ,����'	�HA)J���(�k]��3��/���i ���HI�tGUI��<��f�ϰz�,W�yѣ�x��bΊ��	f����ObPY#8u?s��.�6���J����]�םQ�u�.In�j���F&L�q�)NT�`а��ߩ+��&t�Kдr��(6�ٜ-��O\���E��v�C����sd���V�\���Z�mɦzkK�2���=F0C�r��o��yYj{������ R4KQ��X��n�TG*T�L݄�#��Ȕd����?@M����ӤM�)�І�f�O�����S����r�h"b^�m#�e�<��y}����ጤ�!|h�2�~��s�L�����zM#��J�7�a!W;߭�rCU�T�z㾤y3�e#l"~����ī�I���o���4'ss�=�ϲ����N���ߎ6�s��RX5��e�N7�`n�{S �`m&v���t@*j�40|�F��%c��������g�q�T@��R�<U�퀻����+��q3o���l��2s��#�5�D�$^1cϿ27v�Q���Z �����I�}*���
��l�D�%�P�6���w�F��`�� (�#e��I"L��BP�z���Y��L�FK/��D�C�铝w ��P������YVa�R�e���M��{8��]��ok�/���ج��ԾCR�%P߿��sY�y�X��R���+�̫CW���>�D�"8L6�5å�;�N�k�_g=�x����d<Jx'�R8��cX����0�Z;��]�YE�ӎ�D��7�i���eh.�y����x8�&&�4˙�����D�������p�ouD�>HQݜ���t�#�K�_��Su�Ǵ��0&��~>P��Kb���a2����J��1�V�fc$'w��-�[	�����6�s\��wϘb�-�5���Nf�x�*�q��R��V(ջxrػ�9ٗI�~3L�NoX�a�)�W�K{���}!}�d�	�Ȁ��{ӯ�kJ���Ag���S�O�z�M���Q�۱ȁiw�컖}�kl�^������~�ޤ�A,��BD>y��n� �u�>��wM5y�G�%�|�ce�湡V���vTZ&�wH��A;�퍡.5����,Ǎ���m����ȝN�0N�#��9K����L�	f���V=~<��DQ♴�x6��4(�W�X�H-�� -��k�*���m�3��ÒG�U�ۯ�ͼ��w��EK��ڧ��/Z���p1/9�u�;�p��ߍ��N�G云�]B�l"����m��t��/2$
�����>����vFW�F�cȨ~��Y!Ι\ӂ4ɓ�X���ĳgD�>l&��V��N�HV�j�\�?o��mѿ t��,|�j8�PRH2����ïh��Z0~��'%��)����s����HB�w�ރ�r?e��&�mH����ׇ{�'�ˡ���.l�,'"�D�}��mo�Ͳ�P ������R 1�B�ڀ�CV[��9y�u�f�>�ߞ��w_�N,�^ ڜ��Dq�	�ԃ��4X���p�rѬ�"k=M�f�c^�F��T�ΐ�c�:x<a�,��"`j$#c��Μ�0�WP����9�T~w��P��YR!�����Z5�S;[PF̞+.�"���u
�s�ط
�"�1�X�+#������|i��c��[u4n��Nx��{��tLJT�G�F����h��B)T��ەqY%�j%���о�9�[AM���c�@����'f�͸�a��0�e���5eodۋ��;����"�\p�O���igv�t�h��M���G�t�6�XS�ZQ����@�wXlkVLt��<I��z��)�ɩ�sI2<7D�����d?L����#CI��3����g�o��й~����x�4+�_��`��kT�JF�����%���`�n�%&ZG�"�?W���6U�X�!(���m؎eRf]L�(����r@V��2f�]�+�l��rۍb�0��:h�����n���R{�'����@��K[.��Tc�Z���#%b��n<UxP�Z̸��Z\�`[�W���k��٬��RRJ&�%"R��gju��@��IS�e�Ud��Y�~�zA���D%��$j����'�X�`,>sp��K��}�j�Db��ō�"HY6O��m�T1=Z�������A�Q�İ�o��x�5��?�����&��t:����Ѱ�(��r�C ���7C�����^ 濰�>s��)vU�1���A� #��~�t����N.�@����֟�u�������[H1�v��O���#��i^�Is�� !��6�V�i��?�=�V��]�6�d6����p5���l�Yv�0���c�ȯ������'�S7�Ez���\�\\lK���[��+9TΘ/�<���?"Ns�ݲ=E��E���}�F�V�Hz9N��s��K�0}
�ߨ��R,Z����z
�A��罝v{�>���L�?�n���_ɀz�r�;6�n�P5v��0w��%�#��b���ጻ��8>�9�(O"a���ZfZj��e�'�S�`ּs����y�B%Ҟ�D�n8��"���T�v}Ic��c��ejR���IP�YlΖf+ ����}�f�m�����+J����7Z#&�[0��3�)�g�2����T|�V<�|q}�W2tZ̵�����=�39�߂a��-?(=ʨ��|{��<���4+�<)��}�F�����ϭ�CY��p镂G����\�K��O���>��Q�d;nB�'�1�PuZ4Gw9��[d�8��hM���jC���կI�*L��8�,˵j�i{�9d�ȧ]�Mw�1������؆�OJfn�eF$A9�hpz�ȏ�_wD�� �6i�����9���C�_�/�oƳ�2�� ��K��n��4��Xh�ٻ�z�ڍˋ,��z��"J�n����zϺ��k`�8\���#� �Q�t�v��N� �Bm��`�lE`�����:>3۪).��6v���T�D�Ou!��D銻��e6�
�sSp6�xa5to���.��uh�\��cj�R����:��<B�T�3���kW;o������u���u
��a���g�)��7S3zEDYF�$�����47��G�񍂟�Ri�����F�SQ���h���	�x�h�y�2�����>�	��H,V� /b��P����y ���3�#Ƒ5bDX�/��"x��&��]����'�ֽ��.rn%��q�S0Z;M�Ÿ��Y���+acO���UT![� ��o�0���F�����H���k�o�l���:�@��/�f�Ǫ�}����K� ��:~�4�?���g��ZJw�/sNKr(��t�w�ʽT٩���]eC�ս/�cu��	���� >m�Af4�y�p��b �Ir~��VTM���`3|����S�7@���X�.�}8lp+���j�z.?�,\NS�N�����5�'HJZ��n+\�K�t�/�+���D\�j���)֍t�B��;r�N���_vfl���6M-�N��o���a�!s7���K��׫˾�{c`��^M`zt�h�я@�N��߶\��1>+�x�(����?�2[Չ��c(Eۻ�ZB
E������QO��.z�R6v7��ʅ�Kzث&*ubڲ��ǘؓ���J���J{�l��Y��=Tnh���J���u�<�tr��9��k�ݽ(�-l�1��p���wK��U��ߓ(O�$�/�� k_s��4W�t2xq��������H[��ȷLb��-�Qr�_���&B��b��6�q������i�0c��b�D���^��9�ۣ@n�p�
��ʍe��%�e����h�QZ�_��~�+)+� :.���cU�= Q���b6�#��n ��6�:�L�Dn''af�9�>W��e��+kˉF��}�0Pɩf9�^�:�=H`*T]<�_��%.}u��X���I�b��2(�QTR�C���6[#�!�O�]#�P���U, �*0�|���%ϥ�e�lN.1���lI�Z���Ŀ?�(0��Oes�)>��+]G�&�a�7-�/@�����k+f����2.��V�;�9�/�JT=���OO3���L5Ud/ݺ_u|%౞p�Q���e�g��y�C�aK���g'�]��/�F�>O������@� ��pg/����Ne}.����Ȇ�>����M�����j�שx�ٚ�8��9챓x(�+�T�CC��FU���� �읏7�z������ sJ���w��VC0kwK!�%9�
��׎:{��Y���q�S#��7�����^+�I�}��^^�(�91
M��m@�_�:&�GI��:%V-��NH��F{n7�1 �J������a�ԛV�y.�p�BO���~S{��8�������m���鮚Krr?`�"��;���^zc���<CzK���rjW7_�=ӽW�u_E�1�}��c�>�~���W�l�O�F��8�g� �sL� C䃑�ط�(q�8<l����YH]8/O
-�]��޸�gj�5�k��v�r��?m�&I�U�T~�6�f��7��#�x�B�y�[�	x�Z���Z@Y@���%�J\��O�hJ�/��13q�?j��U���ޅ�Rs� �C��	��ƒ�0�'8�f��j��4`Ņ~�.qB�Wp7'X]�+���l���{��Z�%���A�ڱ�. <�Z����s:���N7BmH��P��v6H�Fx��.aKyp�B-i�<H�C3ItŉA�`a��zn�h��0�9�:8EBM�[S����ms
rh/<���Rg+A���!�?��ʬ�}�gu)�����8���Qa��N-ӊ"F�������V����'�� �vI�1�1��is�^,ӥ�y�"���?�Kq�;�:�:+��j���~��Rp��:*V6��Y�P�:"Q����bj���/�a�mi���J�O�Ye�'�&{ᡦ�2l�	�H�Q$�،#�9%J��H^+H7E�os�a&�\���rv�����h��;�=4�_p�a�uO5��ͿbiA����=����-�V@n"��0ov~\쉬܉y�}DMZ�[��.��E�f��Y���7�T-ˠ<*�5J7���j��M�&-C
	�����2�#q��F��a_ ]��m3ޛ;jY8�H���g$�ʄ2�)���ք��{�3����l�S-/�ht�Et�34��2�����9��֑?Ytn�x*I����G�A�k��b�.�b�a�gޅC
��vR#� ����زdk�:m��HBn�%�G@��aN�?�5��6ù!^�X]/��v�6ܟ�+��yGx�㻎�>ھhf=	݉����<f�-	��'g�tN��'����r.8�\1u�2����d��lL����F����f*x�qK��Ƭ$��������d��)p^��.ʨyf� �ɣ�=� �b=u�H!��y�s�ڵ�����T��{����2�yJ��y�,]�/�1rϠ5;x%��Ya���R�(�u��tk����*�h�&�=bB��gӹ���	GP��I	e�o��ʽ��������ڏ�'�)�X���Z¸;��n��S����I�V5���;�
������,����U��þ�wc06�P*1�>����w&~^����n;������=̨����E��\�t_���U���US�S*��Zz'�걶��i	�#���X�+���8э�m�7`��dɼ���V�la&��a�p������ݐ�3�2Y��+������fEj��1Em��]4�qj�P21��,��t�&i�\6W����]�/!�U��C� å�`�g7�t�2��{��̈���g�%C�e�w���"a��c,a�Hg=!&U��$d���"x�0�� Ht���Q�=R{��	���QԤ��W��	4Q�e�{�����h����u'Q���t�fyE�^���00swt?p�R�`[�^���� �;6�S���l����c䆝��V\�r��h����y����m��5��	FN������k��(-5���Z����m1��b����_���@��>��F'�IF���T! 4'�q����$$�s*M]�Z���s�OF�憻N�<=�ӧ]�%��Q��Z�#�B�C]��>�ٻ3
jZ���'��cz8���c�l�  I-"8؄�d �����:�"�H���X����kH�2~>X���]��~�����v�m�b�E�����(Dt.�N�m�y��+}~v��)�`:1	�U�aE#�3:�xz6Di+S1��"yb�:v����L��Dj�K�KeR�ƲsMMT�[h��}�MJ�[���j��0�@�Ο�"I��_"ύZ.dyP3�E�/t�l�~�5f����i#�0�vX����;���,�x� ��0ʺTv�n��
!h���/��9��[V��w��M`dhї�;������ּ�W���+�o�Z�xP�">�pmC�jc�8.,^H\G�<�i�Uv�w�0JG ǆ����=��0�WI�H�>���=Yim(�/����}9J��Z������ݛ�xA��ߤmkQQ�'�����!uI��i﬉
��Z�%K������z�Sr͐�}��OA�4����(q��J��y[=�K	G�ű"�>����/%�p(qF�����a�j]8�گ���f:n�&�G���e��``cc6�#�Y�IM|`�no��_YAyY�o[��,F
Ƈ�_EN4
q��;�@��>t��ٌG���Qcj.��o�3�WM����`MJ�0�+@ӿ~;����v�8�e�]h�E�E2�U�DQsN�q:������x<³����%@ѓ��3��w	�&�/��/[��-�FM%�(�k5���QT��:����R.��F�2�*K{a�<����#C]�i\Ò�r�q��o����R�[\���m୥�o�4|�;w��%5τ�<�}[	�`N�Y���V�af�����l��>`���I�ݚ�ݸ6)"���Ӥ023!k�B�5�c?t�W�1��$���K�`�'�s�d�K��^���Zu�c"X�=遌<'����ȼ?���ȼ����xRp�o���$��+�u�^<e�r��b�����H\	|��"B��z����0�z��D�$�y{�Q�Rᡍ�L9KYC���<�c;�-^2�m{#����������������>Ǐ%a�K(���b�c0QqK�C�B]c��G`�Q��3��Y�y5T�!>���*��DYS[	�v/8�� �ڇ���$�4�����^�F��3^��gr�:�
�.B@9ıq�����(���Q+o��\I�"6�t�6���Fƨ���dH�_����\��F\���0�7f��c$go�_�#.���8M�1K\y\�[YDi~r��P"Q:2=Ȫ3��zc����d�v�ytaTÂ!���I�x�n%��Ue��aa�6�5�G��ҍȢxM���W2
;e��þ����7��WB~�b^#�S���$P�<��+��}5�r�����ΔE �@>�VY�#����Ba��B�]�/c2�l��k����P~��5�l�2����<����%���1]�[+{�p,�,��Y�*6I90R�(�F�
����!c\�O��u��Zs�$iL�-[�Y����]�Y��j��w�x]9q)!:���mi�r�}đ�l�&+MDh�b�ۻ<��Xŷ`�\W����~M9����w��<M��)|ܣǔ��Yg�	V��*�������K�)������7?�����^jw���L�r0�I
�INz�`��u�|��U�����fز����
�S��������b|�n:��iH����b�p���`n8�������Ꮴ��P��}��M�CM�����+��D��J|�q�k�i6 �mߊ}��8rs��r������+��g���@=",�PD7����)<����N���I�u�U�ݓ�y��"�Q|m������:*�H�s
3��ԧ�!�X����m24�!�����gM�����Wn�c����=�կT(��1Oq�N�",�u�k�9 U�j�D�rR�O�����א���p� I������^x�ݧ#h{s���D�3�=��>�܍�Pߤ2���|y����f�gIt�|�P�=��Z߾i�@�G~�m�I��绹��֍�F�˻Z�	���$�'�,ò��o�����1	��[�S�_�vr�L.0��zZ_G⅏�Y���s<�ɏ&U��z�v�10���B��bp!ר�P ���:)Rr��Ou�k7u�?��ƛ�3��~^�ϔ1M����vE;����^�pw�oh�|�F�Kp���Ц�8����b�!!n�����H����W|% �@����|^����;E��id��0�6[Q�YY��tdP��\0:�h�7����D|>\�v�;��)��^���Z J%U�����J�^����2���TU?FWbZ�]�3�{��貓@����'6��w!�ްj�nݶzX��2�,_xn[�;?!o�M����m_�ԋ�p�~�~(1�'-D.��,�_�v��y�x��o�ʟ�"*��?�8��BHZ��:4˶v��]Ċ__1M��`Y�1���]3X��#=����B��2�N�$VΓ�LW̢�ߥ��8Ԛ�}ֺv/6��(�8Hvܢ�{��T�+R@@�"��4���RV�#�o�~X��1nC �n
Q�A�I4|��p��k�	T@j�>z�2s��� ���e�x����W/�Bp���*�:����|Y[�� �e��`6��Ȯ�t���+`Uy'�����f�[�� ذ���KX]��N��z~�@������[�0��Dˍk���\�����OǓ��]6�0��G��Z�Z���z��
r�Ao��l�.kzeAR0���Zw��K[�����f,�ȃ���A�E�u,�хq�e��d�Y>�q����F[�ZV�
jJ�R��Ы:#EU�n�����K ��-�wC���O;�Z��9 �^�[və��N��ņ�!��S:k/�sN煪�V��Gs7MP�A;T�B�e�J���*�AsW�*o/,��fI��9�9�փ�u{�Xn���)���E�x�`�F$�	YEmԬ�������w�������n�֝1g!s����b�~O��P�GF�/�RuG�W��a 75{Po�?�(2T�����Ν�}���v�+ʣZ����^y��+�T�ޙ�����k�7��	.ڏ�fd.4 �0�gQw�9=O�:��?�������e�l� ���҅t�)�hF��.���kg��D�Q���bN2g]�*��L�C�.�1H�[��ץ�/!5L/o�|�ѳY���",������H�*��*]�ӻ��Z�Z
x;T��%\�*�)��pz��%���=EW�e\nu���眔�1����z}��X�;'�[�k/s�c �U�&���ڶp�NCJ�� $��k�5�Ⱗ �N>��3�w��:A���w�e�@r����?�q�Q���>M�;�b?F�qډY���(i 7���zz��kP�i���u!�,�}��>M	��!���r��m#���as3m�{�a�K	!82L�A�����\������^�V�+`��=�V��P�i�A!����բ䐉��3�r`?	���FBY�vkd k�ѐ݅�ۦnI_�:�k<�}I.�3������O!�R J��ɖa=�v�	u�Q�?�v�N����x��P��;�N�����8�7qȧ��pD:�Է��T�y��}���:�l������N*�G'k�VL1�4z�+�/T��1
���/�;�z"�R*'@��*
�[p8���愻�=�l��%A**e�rp�$��ҋ���u
C~��$nS^t�+w?�`o��v��e�i�Ҵ�Z�0�_n�wpVU�f�N�u�A��51ܸn)&ƒ���y��1�#���A�+�g��RY �7����I�R��ym�#�	�l?,R��]Q7]e���.��&���mH�ά��, ͨ�?��"�>��K'K���/���(@UK�j��|�xRӘ�����+��~V�mp)�x�N���4�����:��,v�	;�@w)~Yc�H͡#n�ZՃ]pa�S�Nn3�JN�^�J����{O�jw��V��l4pa�����0goٌ��E%��	��K/K.]e����`+��s�UČ댐6i��g��ż9
u�Pl�u((-���`�=lzc4��?�W��A�Dޛ%1�F��6#�L�xĢ�	�H��>�E�z�������M� �������� uU�b�!��7�#�v�yO���X�&����繧�v��í\�n�T�ĸ�h�+Lb��l{4��;s�I��W�`#�����1��a�	~B�����Ϭ�r�����:cJ2A��%Ql�� N�kP�!P�����QC'/��G?���-��xML�� �B9��Q�K��JqM�"��Zk�g�ߤ2W�����S4�̼;�F<<�1.&ǅ���c��7�i��bx羓���M�wr+�>``8��󜌪�]r���*�x�_�s?��0|\�=�O��=\�%J6?y���ETsb�6=�md�u2:����	�8�l�FKpJd`:�4�WD�&� �����=k�}���T�
�P��#f�]��@J��*ǧ~�D��>�t<)P8scO��r��EY���ko��t|�'L�i���Zo��]� �P���!���)���?H P��R��}�ؼ�Å����^�����W�i�yG%�/�xP�7���Ǉݜ����!n�e�hU��r����U6J�0�^��*�^�W�4���H���NP�W6VZc���=�E��pU�|+ �:��6��_u0`.=i�I@
OW?IH�(��:5�;�Up!����X�V�U��|�����l$��p�����P��Öͤ����z�G���N������1�� ���jh;N�OQ^���&�. ���C1��[q{`Zas6�"��?w�Nkt/�^87�<a���_$�=o4ο;��<O��}�Y�� �5$�!`������n���isn@|�LΪ�>��認}@��W*|�ad���G%*?dA���|�T��6����/��k�ш�l��fݽ�=OF�LU�sty}�h���f�s#M 9��z	S���NE������ύS�G���E]������ċR����T20� V�jO韮��n����&���kHMܛ[�Y�N�ã�j�~Ax%���}X�]��Xy]E�Ș�Y9V���ھ���`����.�o��%��Ovwz����T�����1��f���d��Cy)�%��P&?nb���\Xq]����ڞr��dt�<�.C6k�^K�jv��,�#���)��q�^�፡��)���� �5�oW�R�(��"�ٲ����	�@��8����	}Yv"+.EK�+j������w���X9��6��!T��ۙ���F����a���՗���r�2&YK�d۲�V��.�'+`��z��4&�
�J&|��w	$)���Y��)����W�P�%�b�}_	��,�[>Qޣ"�Z燃P
gؼ*U�f�eu��4���;i�U:�B���6D3�K�x��h8&ײi6/x�p�ef��7%�,B�I�np<J�2'Y0`��Q?��^��m3��mA�$��G�\�G����7v�|��j�UĶOMovI*������t=,ӟs{.؀�*��"<l+5b��)��A��I1���,0�yuYl<����G����÷ɑ�(���0�O���~���D�L�ë���	u�@u�*�ҩ*5qxn�+(��%bm��窯1�ȼh�vҞ=�)��IX�Ժ�zM%���
�r���ϗ��<�ό�3�	��e\�^��$�u�T"ʧ�������q�9 ;{EYs����t� �h�>'�A��&���O�ҵ0�
2o� ���՞b!{?����l�Z���Q:��ND{?O�|3j�$Ӧ��`0�.�U\F�Ǯ�C���@FJS^�s�_�+r8��>,K�{�ۅ��ϳC����wY�E�B�+�ո&��r��1ʾ
$���`�Ǣu�s�h'k)�����SZ�*sZ7�?E�����O�
�A^o��.�9���?L�B
�_�VZF3�n
�.�v�D�j�D�|ǌ����)~��y>Q�=>y��']fv������ڄ��P#��i�iO����f�Țc��ԗo.�:�9D���F�+UO�J��N�tEz��VfT��D��Ѫ=����fI�h;�l8,~�	�_�fI�CK�;�e�a/ԁ�����V4�i
�)ծ��T2�"�Dw�&a���N�J�a��4��|ׄ���Zka��px����`�Vڥ׽]0Ty��VU�Z%-���%�����kV@�Q����l��
�,Ul:>�u���1�e�1�8�pLpA�SA�����Q�i���8���c����ۙH�^���ؕ͗sD�g�W��\�lO�E�I�7�3��i'Y���ͲG���RN��ˀ�+FL�]�B����J	T����뻐m�$%��|� ���q]n"��Dw� ��Z[�`3���,"�Q��}*I�w~~��1���s
`K�F7=��y_�&��kf�C����V@��^��)� �I�N"x(d
�ˤ��70i�՝E�σ\�8�Ǽ6uÀp�y�^��|��z·�%+Y����g&�g꽹ҳj���������/���K�]�b�W�+l"�V�ڙ}lc��K��폻�Y)���S߽ʟ�Y���;}�FA�2Vmz��1g�dz�|
���^���b�x!A���xnu������r�6��[�����d��Dg/�o�d%֠#�Q�ݎ�Ԅ"4iD��f�JEs?�v����w��}y���;�q�"�{s#b*� 	�웈����0�Ոs�'	�T�i�=�!�{u>ě�g���"��0�e�.@W5��n%Ѱ!tp�o��t[O#�Wo���~�wt�-�б�D �@���H8��݈44�ټ�1H���o�Z0��Pt3�|B�ݹs��Q��Y�y���������8��Y���{��be?}�∄#]uġw"��+Pz�!��Q�m����^�ˤ{����Ϥ-�<ľ�~d="Ķ�󐛨��M�=u�O^~�F�N�t��Ň��e�g�4�P�eYb�C��=���c�6���08l��б��%ІQ!A�5oC�}.���Qj�C�����@<�!�x�[�y4o7T8�/ ��S�
G�����H���^N�}�ӦY��Z+31w���fˀ�f	(7;�v�������@~��Ǵ��Kύ�mv1��T��n)"ij��
���C��ڊ����q���Y����O�@vOi|����="�w����Vl�x�U�D�����┰�i�t�u���k-L8"�D�UG�j���T�Hm����l�sb����!��e�&��d^�-�1��o���>�eoE�=g1��|~�4�UE�E�u՚W|N����9[}8˛�,��`X��^�6G��ɹ���iEsl��4��+��S��ݙ��,�X��|���R�bf�Wv���V�+�IA���w�C?hd��u�~��L����t��ל�;l&�R�y:��ع<�B�=���CAv<��xDސN�xF[!�% 2��7<���x�1J���%A��)
��Ƈ��biZ���&^..�Dzd����u�հ�/t$|y%��e���=b�<%	�L���\��c�{��_�v��ݽ
��A����-w��ĮH�w�W�0=j89�F�$9�UT�c���ب��&�J��ąixV6%�5�:�b�mQ���L�+��Xm�H��Vfh�b�&║蛩w�`}.����5�Cw󳍷�x42f�&h,�F��{�y���2�4%��e�Z ���m�+��li���[U�*�A��>c��
�e9M����'�D8��+�/�cI�w�q��EHj����7�$���$�
��4��%�Ӝ� 2}�>6Z�O�_u_Ҋ���׍)HF�L?� 3�:�����mk��n5İ�el
���T��+풻/��Q�@���4QbcS���+J�F��; �)3��5���7ء8sQ=Vpf��������`΀�Ku�57��}��v;�nCM�3��[x;i�ྫྷ�zN���#C�t��Vq������}&�d�']�� 5�oUh�:_��(�v&:�Ζ
L��}w�Y�[�Kv�M�M�_ZA�#�kUQR��t��8���>	b����.w��^9��������<"�B�C�x��y����x	a_�,=�x�Q��Ƭ��O4�H{]2w�}���6�m*�<��U��`A��x�A��3���j��s*�p(B��X�ޡ��W��y0��4�'h�����O��M���+Q����lbm�q��zyq^��J���h����7��gy6r'��(I�d��f���2A��	���O�r��58�'O^:����Sj���gr���T��	�}Ӧ,�M� I�d6u_����aZ���S)�.�%u���:S�1���z�� �*�i�lR��qQ-���Y���8��pP�8���Ʋ�ݝ-,.�p�΁P0��ű8-G��s������د��꜐K׏y���"���Z�O<��^��X��\@�DH{����,�]B)�`G0��;�3�X��j�Q���c@C,�&ज�6�J�Ad�:-�2n���NB�o?���@�9��W�`y���-Y���,�J�U���v��d�u8|���3�����
��,��y��Ŵ�8n�M|�B�r�����QC?��>D��=w�b{���7������������V�Q�j�Sg?6'W���#�����i- 7p�?�"�%�N���X*�/3$��ID�yr��-q�MțD��s���2��Ѱ]�����Q$~cD�Fo\u���I=��<t}�q�6���$�c�V :�eӀ��?�Fy���T�bU�BZ���t����Yr���èБ|3щ8J�Xd��Ў	�p���^�34'�F�� ֫Q���������|���ҫx~ʁ�m����"�$ϋu0�k]����6�� s���MF�z��$;թS4X�sw��`O-���\Jͮv;��E�,�嚹��?~�c����EIm?L�~���k�t�}���a2}t�PC��2�*��/%�dM2�,�ڿ������_;%$;A�{A�O׬���Ճ������6v���Z����C�qD�մ�k���m)uL(����IJg�﬈�6�J��"�A�F*�r|S)Vm���N�3[��2Ԙ�	�[r�zD��\?�8n���f��<O����<(�����Fa$��s��FM�z�3���!nyn��������c �^Qו��V���3K|�I���m��wH5`k�f�~y�d����RF\�R}�6i�U�?;7Wpk2�u:��_-�摪7=H!9�P[x�:�G�MR��L��)����q}1��e���S��CL#�����!�2�q�w5͛^>%p ��t����3��j��}��/$����{�ʷ }T����EX[��#��K�|A�n;%��~�5�/b!���
�yWˤ��fr��:����3>S#�t����"��&�M5����d�T�5�ĭW5���XAo:��4��9�ۦV:s���$B�HF�um��n;��ԡ�\G]l�XP�B���]zvzRL����g�������s�?B�Kz��w����( G�'����7�.�Ms��he�����)�=S�0	��s�i�.�:h�/uI���˜O8O���vt��|Jn�jcW�F�ZO(�lӣ������z^��&hC�Abb������˅�#�Ȱ�R[ީfU�ii+�៤�:X�:��۸�F+�9���Z��|�	�����G˾��ħ����:�pO}���/a��R���ܯ䣞��¹�'�+��8-x7��=���s��XuV���_�z����q�5��'6	��.�ܽ�'[�d;��ݏL�X�C5,^t�Fb[n4�n} �~)�
��|P�~%	
U(�ʋL�pՃ8G�%���ǨP�[oO�F'qJ-ZoU�OR���L��-�V8wA�vlJ$:��]�p�^t2�?8�l�ot�8�����S�ńgOI�K-y.�.9����$��	�`�����B��� c��� ��]�2�����&(?�}����:{�V}�9����������.U�����n�ua����0(�43��FnI:�<H��OR�A[V��b.��^$2sF�d������{��mP�"B?#5zTC�
��_�Ť�bN|xO� ߯-ŵ8��N(o�����F�s�U���w��'�=�	�=P��g
�ʾt�I$��aD	�7cN�4{�vƨ�Q�ȗ���ũ����&��teGr��e r)&l��R$c �7)� g���2D\0����N�^�������y����p{��D2�p���]t.�OQv��}~�|���`*�5`WQW����x�K�r1	�c�.�\�����p�Qm�]T&����[��k���)�'���$Yg�P��Gp
��W&��Pʽu����fZ�MN?E*	�6tٵ��J������[����)Q��\t��y��/��xʆ�{f{3���I\'�lɘ��"}�"��R�Ņ���<>�]��Q�����w'֩��]�JT����m�U�~��0�6,�)\�9�v1+��tZ�`�q��y�1&�n%�g#�^�≶��#�|�f���?����+��vn�[{�����`�dh��tXD� 9>`%3�Z�Pjt�������Ԅ4�]}�M>V<S�[�� 8!������m� @��;8��S�N��k^��r�y�&P�A���t-ŦR[�U���#F�Q�Tp���*�����a��8�D}�l��}µ?�:�H�j\<��6j��������_/�W����Aӣ�g"d���#l�Ep)ʫ�(�4�ElQ0y����%a^��	���i�S{�W��tJ�<������i��v��O�kO�<���	��4�%����2�H	���Cԗ�����"�^�Šz�F@IJ�ć Ӈ��U�0�M����b���G��"Τu�F����b��Y�j�gK����v���
D5��P�=�BzZe�CF��%�aS'���I���w�v#ڬ��. ��F]r�_K�����8�Y����j�J����Ck@�[�P�.��OǗ��P��4mt�� ϕ���'����LHa�>����n�F]��Ha��%=����H��:%�U/�
{�%_� Mǟ�S�<C����	�^�)m�� Caګ�Y���}d��)Y7���>�J�3�L���jQ����J��FeK��pw�9�aY
�"Ŵ6 D#- ���#��μ}:Йf��L�c�6�Lh�Ya�*ޑs�y>`j�uN��2:����J���!�ϙ��x�		t�:������K��p>��n�e��i�B� �u���,���Z!���qѣ�����|����s�=J)d X	S��Ui����U�6�:1�n�z���$�,0���~}>��u�Ec9�a�j+N��#��)D?vI��x�ǠШ�ΐ�D2�]l��R1y�]�d�ê��O��B��f4{�K��[����[�m�B*z��y�W��[H���M��i��b��e��+��1.���~�rR���!L��cz��>w���D����~��&--V�
P!t���+oȲ����� 7��W�V8F;R�5��O���5r-�W6];A��w����xω3ǳ�f@�i��A�暅)����8�c[���ͼ���q��[kq?_dyQ����`4�iA��o���p���m� hf �� G���*�4�M�j0�׳�9M�|,x��bA�'�+4zcE;.�<�@��
��̟��y�>��#�{3��[��yI;;I�������MM&5?/J�9�M�YL���Ϳ�b�a�Є8I��9����g���R�_�ґs��t�h��x�0����֐��f4� a0f�sˡ��P�S�d��#��#��q��=؋����e< �Y���MG}-QЦμ��)�����t�&�v#yDV�ȐlI�
c�@���,(��B~�h�OvpA�B&b�W������`��S;�夿�/t����mbg�
��;��5���c��ۀV+X�(�)[Y���w�t5.)�/��g<m�ꝵbbX�2���G�R�o�_���M���	r�zs������xw��)�j�ç���B�̬���i �D�K��8���>K\�5>�fQ�]�~�+�+G����~/�zsB�������EM�^ߩb��pFKtSw�Ϸ�@Tt�Of�#ɞ��`�2��U��c���|�������	�L��^Ԫa��%3���=1�_H���Q�~�6�l� dȊ�G` �j$zRΣs��i�,�0�f��S�]�޶�h��$-�7��!3�'l��:�@m1�)E_wP�CU����3֓؛�W��F$��i�^l��iy0{|~�h�G+xޯխ<�
̈́G�#{�c\��#kAϔ���<6OYZ�0_�QIBm���3�&�Y�B}c�@m��iU�z�q�u�Z@\C���M&Ɠ%9� �T�є��%fY�ݫ咍jM˂���Př��{5�tF$~σS�d�����~��%L1�����tiĿz����$�N��h�4�8�6���~�II&{�Op���=�hs%ؐ���I'�"����'����� �'�H��{�:e|�_;�Ĭ�$�c��t�s�h0l�-��+��4#͈�%ȧt�qXR׻�!�T t��F���aА4�#D3E/���0�;Z��rb?B�x��%��
�N�[�aP��C��#�g|T�#{��r�:C]΍)�t��Z���/x�V#�K�������Ŧ�`VY(��7��J� �p;!z��D=�J�� � ���e�D%���J�_T��"A����>�<� �5���nD�皅����l�B7IC6[�ÄQ���֏{e�
 ��|�������k6��1���nբ�8|��ɪ�@�!K�@W�Y'5@I�鼴VcU�y�0C)�hG)`�>����f3�+�{?<�é�e-�A��Q��J��cdm��8�?��2�{׸(�MEH�
|�3Q[�����D�/8?��kV�6k���
B�~hc���d(���m�KѲ��5zۨ�k�,��2����2�h�Կ;u����X���{߾��X(��pT��_J��F=��#�`���'�7e���a���3*E�����m��{��4ƍ���t�D�r~^ E~�#DT����� ��ъ"��gǠR�A���"�J���e�9��{)�)_*/�?4ц(�Qj\�T����S�a8�+�@���S�
�?l�X[�[�����&��u�50��&���9wa܍�,�YN��D���oY�J�J�9]�3�-�h�8��U�g����w�lRSP�׾n�@�h�O!���7���v���B�q\}P{�7& ��>�@W�@�� �p�l��%�R�Ժ�l8�mp�i���� ci��5���񣺓/��<|�	��?��
�j��}��ɏ2N>RE�ΐ6h�m��U��n����ߤ�N�Q�Ы��i�����0�l�<��n��Vd��h�)fA�\�C���#@����b���&�l�0VQ� �������'b��U«���b@����?j��=���B�z}he���RO. �׌�h���EC��^O<68���b��ó+TE��VRa'�PLc}ŏ֌8M���X�0�;6E���I[b�Wt�*'�˚U�e�+�� �ԅM(�(�ꄶc�/ȟ2kk_�ܭ~�!�r�,N�ʕ�ÍZ����D$2M�s�X��O�b�p70�[n�O>�J��&��Z `�Z���D�Y:m����4�YlNK���˯�eG�ݣ���(�D�\Q���^� �����S;�/��ŏ/=-��k���S�vw�X���,�X���aǇ�җ��c�&s�&�"�O��#��r<B���?[8�U,�y��~fr2E�-3����dl���ɤΦO{��$:�cmP ;F|��Kk���b&V��n���n�r�P�h�^�%�g����_}2���ŚJl{�ْ�b�go�V/-��mcV��'���"�CvK�Q�^���ژ�T�V��᠖!�j!o�@D9ҏ�1m�����Aq�9���7?bGckZ'�Y �?��+s���Y;c���/��Э+���vPW��mG�*ڵ�|����u+
�����iv
/=�^�e?���~������N��S�rnAi�
�O�1����j�%7�3�|����@�cҊH��eB���R��D{�^��7X��uF��˕�nS��%�'�R�%�����S�q�<�MP�z9�\)���a91�Yt�3[� �`�'"H��,"liH���c��euE�c�{��RL����%�0�p�&�2\F)�|��]	] ���|F��{,5p��c�q�OeBc��́X X�~�@�uU�vx����p�jo:�L.�/�{0]Z2љ��2�Nq�n����t����<#g�T�..��x��C�4�jS_���ס�{
]+r�l0x���s�׆�9Su��>M�n�P˯i��3�P��p�j�L6���=[+�1�X�i�іx��v����⣔�;�#�hUHb��V�����U�&�M=��pN���,!F����#��W9���l?ϰ���G#��v�F ��]1� )F�>��<FT]h��4���n�� *ࠑEG��t��eǈ�v1�IΗQN����=L�� �Z�@C�2j%f�Â
_�&�NF��I���;�f�DD�H��뀼2)@���l�������$�S�B!�P���������d�����������CY]�^ �b��2_@��n���X�\�A�z���ٗ����čR�y��N�	fr�R��f�$m|@y��qܺ�fΙƶ8���
�B\�)q�f�Dk>"��;���ްiá	wM\Su�������u�~o�Z^ؾ0C8�-|*XVB�Gv����i�%��'E���4y�,�j~�W8S��Tha#N�B���d�=F#��/��@ʢ�crn} ����@l�T��E��縴����Ks�X����M� ��6{����r����,T����6@�҂:��zI���^.���r֥����i��+�2�Z�W�s(/;�X5���x�Q�6������r��|g^�r
�m�2F������7�㿾���^�.��ӛ�rv:�1mp��TE��=�eQd}y{�[�i�ޯ	7OAW&�VƢQy������y�DC����6��lG���@�[l� і��ny�`x,�o�5���9�-��v?ڵ"DO*��< ,�(5/�t�вkB>���,�PC�y�L��{�~M��Rg*-�%0a�v¤��0�2�&�w@�NE���=�M�2g�i'	��B\�#��\ /��l]�kP˓I����4��j[����u�$*J��jkr��w�%{?��