��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ���\::��_5x'�o<N+H��}��]�����T*�7������Mk��W�͍:E���$?�yk�46�=�a�� ~4�	�҂�&�tC���5�U�Ht҇E6�\��-��2u��@�d����mw����ۜ/kR�2eX���nY�~1�I,L�&J�B.?��E��:az8o�m�ߩ�M�Z�<����K9Y�j��7��G�o�%	��u~%�xZ9������S|FSFxRO�5}�c�Sy �q2į!�$���<��p�'=*Ҡ.p�M*�\�0῕^�<�A�	��/	Լ"7�5����4ݒ�°w)MoЛ��7�[*(�E�P���o�I0��ೂ���KVךT�b����]:�[��:�4?g0jݡA�My{}��Ǌ0y�#O�H���3B�ӣ~��(;)2HAvY��ն��ДZ��LA�Fð���`��p0[\P�]�t$�E�9?
r7Z�2��s�������K��Gֱ�+����3��Z�s��5��엖�s�.mM)�����Z�6�q0�c�s�:�Y�׽��	g!!�=pcBʖDyl�͆c��f�w<1�9���;�}H.�;A�����M��Cw��nl���d�齤fTi�b!���j��N��Fu��i�~�ܥW���D�n���������Σw���������)�f���m�6���>�;	ЃE����0h,�R
V� T�Y����mכ
�e&pr]o�>��};S�V��e��h^¶���7ߎ�X9�H��곘Z��ְ����b�m�ob��S�H#ޖ��ձ�^� /��
��.���MהZ����&/k��e�{|��=�L $�����>.M�\�Bi�����s�71�-G�x�J]tţ� g93���u���h.0p�PҤNj��	�%�ac#����*a�q	͟Ilº��������HI���_���h��j�d/�ƯD#m��1�i��^��-H6-��B��cT��n�F�礮Q���)»��Z���x��t�vxr4�yE�� }AF"�^JO �p�͑ۜ�-��$ӯ��7� �����#U��*p�~ddW�����5�}��l�la�!4��
��{�i/��?p��P_��P��K���7 S�N�
ʫ4�ri%ф�¹R؎f�m`5�e\r#"��ʐ�*���a����-�'H��Mr�<����6������T�Ld��F?����2�U�x~	�d�eJm�+����;�"���3cؠ=Wr����r�K֎
k���U��Gp~)R�[	��鈂	kT��J'*�	5�_��LhC�(~�=�� �������%�;����O7d�t�����k$5$���Zya uEz���|0L��Nx�Nպ���(ު� ���zv��S�47�tG����W{�ӸM�_=�_*{m�p�U�c̼TH���|���Z��f��gT�6J�%k���#�Jygh#����Ѫ�ͽ�Y�P)S&LM�n=�j�oDh��Ve ���$&���V9J_�����y�|$��kS�c���ҥ�����.����2JkQ3�(o�yc8$Z���Jq���l��Si��z=p����p&�t"���jΩ�W������N�J��}�[�;�qc�\���' �/��|?h�ե�%�#5� ��P���՛L�Voz剩�N�F��f�:�O���N#e�>T�H�)�tڃ;��J;���PG���	$*��S ����k= ���(��v yL|��2�Fk B�Ȓ�	.�D��Ƽ��_D
6ve�U����|�	8��p::��ݑI�9���Ԝ�j�����ڣ���XX�+ ��Č�I����� w��A`o� ��|%�A�C)*�f��J~r�f}�Ԑ2m(�<�Ma2
x���e�(u�*~,�. =�>g��(�}�-�EMC���aD.:�;2�0,$�#m����FpD�u ط(��>�D�[���ߊAW�0��U��^�h���J^@/:Zd��,��J�$�("FXH���+I�mV�?��3w�K�p���I���.�Ԁ�V�ҸxLH�%q�{11&{�ZM�v^�v(tm?"��NFֻ J�NU3��	�ז�fS�S��B�:�M� �w���`��}+��Y8��c�z6�C^����쎜��_�
�"��c�,(M�)��H��D���֗�7P�Y5Ԗ�Z��;A!$��w�w<�JiF$���p��d�!����Ad�H
$��~�]�U��]���[ U���eֿ<�%Tx���j�7/|����>CG��<����CϹ��\"�L����,9@��-��D+Η�tG�e�"x��0�$��\67������������eM�m���!$�������i-�ْ�w(�����M��]LD����M��G��ܸ=*,>�2��;0c�ɱ������`�������/ʎ��v�lhХ����d@7���+.c�3�1u0ä�%L�� J4[�@B`+"��dV��h��y�C��v@z{n�򬟥�)��A����U0^ ���hG������}��Ȫd*r�.-��Y��	����֥j��pyY�7���B욟��AkJ�C��e�
�G�lyV�d?������N�A:bT���D��5���z��e(���K���G��`�9����"7�����S���L�߹��o�2k�n�#-}ꫭɈ*������c���*�@*ߝG>�f�J(���U��ZB?����E�`�&Ch��)FFHR�C[�1���Kvg��*��E7�~�_�t�_ͤ�S~�+N�!�V_U��K���*ho��Mw�$߅�{����5�#NB���hc�S�Cym[�c���Ac�$e�b��}�Cּ�:�2���~��@�sNסO�1�s�xw`P�!�a�+JKc�O�1$Ijֿ���S�ᒚ͌X۰�a��W���O�c�eg� 7@�cc������?�ۑ�g�F�Wu%9Xz�v��b�B�*�$"0:y�9�sïJR~-��\;�i$	�S��h�79R�����bzP�o��`�ܕ��F�"c#	wLM�y1~��?�E��%A�n���C,[�ؾ.�����4ПVX��)hX�a%��BXe^8Ɨ.�y�%"� S������W%Nt���(�j�NN���e���"�t�vz��~:Z˞r%��|l�;;��XV�^^ˀP=�NznNyU�4��i ���L:�Ū9�����#��]��z�GѬxԼ��$.d�՝�y�5/&ů��7�D�;����c>q��1��,1�4���0M�
���A ן�MŰ��7�͓�K�+�-��>��3uL�*vϨ��a�`@�a�5��	��2������=�v���/'J�n�x��p9e�~ǲJo�ZH�W[�ߪ]�b����( �Q/ģ=�����x+T#�`v�I��Q+�RD��ܩ�O�|�h�[��h�F7��A�9ц��q"�$�{ӵ9��L�Z�W��j����=�xNy2`fP�"`��J%��������bc~���r{�Mk�9OjZ�(�:����q�|���)3i)*������ͷ�K#t�ݯ���O��JO�."�B~����-��V�!����!�ҲE�n��!� '�C$CU��%ޯ��}TW�$���"q��+M=��Y�%O}������a�M�ܹ~�c�4^F�o�YCP,B-W|NNGFΩΜ�D�eF�C{y���Ӏ0P*�(� "�;�#��ek_�d��X�"��@%P�C�c4J7��kY!���U[�;?$�w��(Ż6)F���7�F<�D�_�Z \�=.(ߣ��rL�B�S�X����&k�v��+*.8y^2A�=��%��eo㬩q�2A�����NJ��a���eb���֒�
�:hxo��u:�лs�����{���?G	�xa���A���/�{~X���)̷8,��(=E�8vT	��1)�ʲ�S��_�P1���gߡ�fm�ˬ�M���d�x��s$d�j�91�|�n���-�SX~����0
J��r��C62��9��N��W�I=�������}�Y�9�w�x��y �g��������z?Q�Ik�5q%���Ɏ���У���SEuD�:�=։/y{u/ ����P&��N�Yh�����7�f)%1�U�JQ�H���#݅��v���?澟��9��d��}�l$+�>>ˉ�Ƈ��7�1b�/�J=Mr���A���]���6�k��� ��h8?^���������;�p�I~�<�T9p"I�(MA����[�"�E��6� ���M$��K���Gu�Rg�
-��[t����O����Z�;
J�Lk:��if��R 7�\��jL�2���I�Z�>̗)c5!�D
_��x���^�	���oX�U`��n�T�K�Kձ�L��Z�a_�����N�D�t��2�<H��;`�x��+���	�Z;~��9y���E�~�!@.x<�X�?��j�^?��k�`ח~R���y��W99= S5���ЦH�#�4��-.f�A!Lܣ�a��]��~ ���E��A���=�T�+ޛ����-�^��:<�g�B`���E�����H	����Y��b������GiӴ��&1�Q�tu��6�����NX诖 �^���r��YY8�>okղ��j8S8pq��Uۯ/���*}k��	N�����*Uxs�*VD�/��v�v��bg�B|�W����4�l��e���q����O�����-�얀�7[Z������k_t��� �mqa;�>(1.����<��յ@N_��x�0�#�e��{aN)WԘ!����S���o��"<�r\���$�'�=̛Ђ5���o���\j�@u���u�j�0:n�B ��M�l^�e���̞�["���\���˳�+���%�r�j�u8��a9>�5a�F�� ]�-M�V��Tֿ�w�s�:P��F��v%`

8Ѓ*��Zuζ�t�K:EӠ�1%v��;e@K��!�b&%Թ��|*��Nz��~�wDT��2�]���PI@&�wx������=SM�<�_��_yN��#Φ��S���6��*�ƪG�VC�� ��&��+O�q�	����a�r�ZxA�uR&B�8���v,V^�ۄ�m1��̲X��%+p���#j^�0j��^(
�!��nS%Dc�wj�	u��/[M�7uH�TK�]�[s�<���~D�F藈��Q��,���I'j۬�{�w⅕N�7��1N���K�����k�;���c���qA���!�����m3�$�Z�k~7�4p��z#u��� s�,�A[��pQ3��+���a�myP.$�yK�Q�l�A����eq~Ę~v���a�U���\�J�3K�0�����;P��{u�^E\������M����觥����Rd�u1e!���P����ѳc��,��l�#���*d&:
J�Q���M�"���rW���
���HAM(@�%����2�3*�w�>¦�dR�Y�=��R*\(/2����zE$X��S�h<	V��0O��e�Jf�dK��C-rY����	(�p��z���<&�]P�.fd�r|�=�_�\ҧgI��同`F`X�7�'�+�xE�]����L4$�*��7-��Z]n(�,.3=��(�v�t��[�0��'���қ@\;��_ ����[ШCﴀt��VIx�A��F};?�{6�w>�d>k��e�9�g͆b�U�n�S�sF
�=6�6�.`��l�j1�Y Ic����:B���r.|;�a#劭�qqY95o�_�P���e�˝���v�6��E	���N�k�����z��
 �Xŕ���]�*;>Ɏg`��f�j������*/=�xr\#ײr皣!{����SaȒB�,߰4��vJ����,HC���gW�E%�+����͘-�'_y�85�J���-���VH���R )�N���#�[����7_�?l�����m㭥���ߋ��`u!�T	~}�[Sl�������:�DȆ��z8P���CP,�6*��H�*{ڰ9��&�՝�c	�
dʸ��/D?��#�v�	 =��+��a��8Q3P��R�
�����;w}��'��%1��w��=�>d{�̬X��ކ\FK�!�o!yP�����b,X�+p�-���f�R�F�&U�߉
�`�l1+�}ԱM���H�_������\�������\8��b!��%�ycD�xG�F�f�YI�ފ�����+��,L'��*!>'��Ҵ��F����R梚`���8����Zr��������pB�c�v��]:���~h����é���d��N��7r�����^<9@R�JD
UT��\j��o���B��V��:#���'�G0���?Q��JQ���j�ݺ����X�L��M|���ob�ZOم�PK�5�4�>�ڃ�ɀ���-��¿�d��y�2w�U���GϢ�Z�����,0I�� �,���x�5��~����u(�l���%n��sqO�[򏳵=0�k/�mY�-P)�����E$y -.�$�g�A�����7T����t�9��\��,���d�6� Uֻ�$�^>NR���c&_3YA10���k���Gfm�г��Q����S�=�#%�ٱ��BK�b�X�
��B.�@l�Y�: 0��X]}ʿ%n�0_DV�4��mED�'����x/0-�����n3y�Z�I���{~h?ܗes :��=�`��W: ~��r��y_�<$`�P[���9s�����65^�^7��M�s��Í�L���"�AμqxZ�ԣ�* v��-�q�y��Dt⽖��=J�'���{x0`�Y��P������0K����U��e6�'P1@q����'-��x:�@�Á3������,�������3p{MH�v��\����;�<K�9(���W��v^ˣD��琨�|<���M&w2�*~6P�M�v׶�5j�8��bZ�Ƞ�(Hfw��L����S���F3,6wXҊ��b��o֎�Q�R;��������
�b����0���n3Z
����&�����{X����[n�p��^5��*:y�8BkI(i�n����ř��lR�L=�'zu1�4�6�YZJ�R�]���*<���)܊���R�t���w}�5a�@��6�'7��H/������5�d��iy��81�E���'��Jׄ�^�A����2��������t =k�FA䯣���B��j�4�^��n��-�Du����4�I�J-N�Ci��M�?q �mm��G�ל�,���X�Vt��n2�[��`�������x&7-���y�Qp�(U���rŹ�3gU�7ҫ��_ш�1�q��$��9��i"�@uܣǸ���P���}����o�{�ARtk��9�_�M��̼a��I�F93v��aX��92ճnM�d�6^���p���E�r=�ڷ��LqEFpnOb`�%�n5}/�;!����/�2�glRp�|:w-�>��%����ǩM�z�V��z��&:��t8e��WcP5[41X�![X��ׁ^Ql�J
�w�?6��4�^����u�1!�a���G����f��"Ҝ*�Ł��(�nӉ縩�*R��a9����^�ğXa�X
z��5��<���⓿�������W��=|�UK�@`=S\��2{c\EOuby���fgz��v��֒���o��s�_BUBm'T2�YM��{?b���I��.����W<�]����T"5
�4�]ר���� ү�!졭 ��(43�^�:rV~���))|)�?���X?���k>�X���t�(�7����κ,&u���H�X^���ǘTLO�� �<��ސ��;�b����ۜS#��2��a������σ�A�I���t�y����-vT�8�!˜�Si3�|��҂���kCM������Y�����f?�����')~�(^�@���{]��i6��ԇ���nϣB����г`���W�����P�b��"Y�Xn�t1��Mv-����J]�H�<�������zJ�n�Wp_�t�NP�'v�+ ��ڛ*ܸ��6��t�k���碲~"�]4�[Ռlh�y�q������ۧ�S�]��ե��{��
:���
�S��b��E��]Y��ub��8��Ϯ����?�|~^��b�OL,���7A_��`gN�qI���1�����k�|�'�.��99��P)� ?���it����Gv6Tk�f9��,�%�Ofa�Or�J�l��7����$&%V�,�ȭ v(�����fCU�^e�7P�V�ò�B�:�{�c��-�u1y%��#u�W�(����`oZ����U��D�+~�;��F�Mc���;>�J��(Pu�N�����)s?(Ӑ�S�o�a���+���S�r<i��q�FhC�v�rF�5�����e[S�GO�8+��-���w���X[�����7-$�I�21�����65 `��8�����=�')�;v�#�K6K2��[o(�t=�aY�����u��8�
fg�V����kw�Dz%q���\)���n�i��m��KfK�������&�#��}R���%�\�1Dj��"��yG r	���Z׫��"T48��sW��rl��gCX��V0|ǂ$"�< �7k"|��|TMZ��k�z�	�[��TI%�@JÍ����f�w��^�ǫlꇢ.��[wH�g ��#MA�;�@MŢn�LF�HB�'�[zַ���)R�Y����n�T�L �m�$>����N��(tf��J�ІE}�Q��T~0v.B>GS��\���eC2�rάX�*�`Z��Sf�����PzN�SL�0ɔ�N)X�����𔬃)Uw!j4A��g&?U��go����}�^~�����/3� x�$-Pn�?7������<A��/5B�2�v��/9vJ�q���d��_���9��)`ee"v��W,Ar璗T���%l���z���i��Y���
�#��X�����Ut�g��� ��K]�z�^��L�iS���t�'C����cEu&�F���b+N���i��Fy�`�
y���ԋ"Ro.�g?���q$�&��A�ƚ]uaݙ��>Z����l�7�Ӑ��"mrb�.P��T����ż�i�KR�z���"�&�6d6e���T���.�lI��_�m@����؈i�H0D�_+鍠��n55�Zq�yt��IVM���uܿ�'�3�3�ȾE��ؔ?��)�YP>r�w#v�2A���:�lS:��P�Y;+�9-�3�N��D̅�(��+Q77!��6g�[��b�o��˜A*��'DW��c��]S���g�2�m�xa�Y�]����IȒ!
����� X��֒ѱ�-�]:�l���M����,TE��q.��A�r�+7}r�ɻY9�#��T)T.i5������6n���4�]�ГȀt�<7����!a���l�C����	tɷ�+��x}�&
�3o1`��Y��vP� ]���
`�v�O.�.�L|1�WR����{Y�N�	>mS���Z�� ��7��x�G��52ژalۮ�"��ŵ_�������޲Z��L#��貃�
�(,:(��ƅ�'f�J�CBɣv���ӥ�g b؈�&��oNs�{��s;h��Up�Td"D\6���p���k�t�X��&�r�ðT>m���\2�5!�0�f=?��1�I����1��ew"8�k�W5�]W(���c���rA4��3	᫵?�k�qې�������5�M���]��>p�=ֱ.��]�; ��8>5|P�1�N쓦�����d֮9v(��::L�p,i�SO��c�a����qC,�E9�A��f����lw��&TƂ�oh͊a�`��*��w(�uR|�e;��B�uRP�%ϟŪ�c�34���頃���'�Pz ���^ك�E�s9������b>4����&C'V����CP> �H�mư�k��.�]7��Ի7�5Rr����\=M��K�¨N2G �0,��"��g@@��C	�U�h}G�'�ݺRi�d�f���Xeu���9�nA�wҶ'OԕI=4'��_��"�NK�s6b�b0j��\�P^Qj���K��W���OǾ�#%"��q��$h�X�g�+ą�`�3Vx�����@��8H�������$��*���'��p��d)~{�[_�Ѯ&nk�T���PX Sf�8�R�!Q]Wt���D���!����b�����+V͞���i�.�h)zE����"L|�5��I��%���X� �m���Zt5%3�\��
����^�H5�h�x(��"�w������j�8�ֺʜj�� �pz"��j�1,s��[n0׸k�C%bt�vdT�/�7�~

m�L�L�f��[;I�07� �p�T�@�'���M�P��=���@r$��@M;�^^�;l�/�.�̆��u����}v��ѻ�U�xYVCIL��A��UrY�ß�8`�ӫh�p��s�n]�l�eqB�#�H�о�3ҧ���Ar�_��,%|���*�W����8�uݭ�������0�h��U�я[2�qp͡�n=�����~�ܴ���{�Q��O9mxn~�ϸ|z�W�T�k��B��󏥐����]��պ���o�^��P�w����<N�[���]0���ԥ�8�sC��v�3��U;>��&�z�ZʃU$~Q������]����mi�n��d�v� (_��[O����ii��D0ˁ'Usm�֞\+|����iT#��Fx�̜��aU�ݽC��<����ܓ\#e�'َ��$�W��"�u�@_��|��ُ��n�),gx����E���O�K�_|1��RځK%��~EǄ2� ��0w�׷�똡�$ur�g5�^��$�+�W�r��D��ldn���i/O\���b���isO���g.��įvN-� AwK%ڵ[�2mWQ�Қ�9TvՏf��'S�������
,�5�)xa�t�O�Bw-���������.�V���i�c�<i��`1W�^`�g����S��d��-�� ���f��$�sɧ[�ر�Ԃ����%P�U��w�nn(�K J�&�T�>i����c��0q�>і["��F}uR�6�Y�Ih<�N"E���;t%�c�3��3���M����ˡi���[JCOƢ45-h�Y?�-�<��17=�I��^X���2��ooDZ=��޺����m���Ns�+��S�y�,��xط$K{"!�E@۠B7��S�͍�F9�� ԥr�Er���Ya�f�7�=qC�֋u->��Y�~1�]'l)-�}$�ؿr���T�x�1�+W�A�fcX.������P<���.����&�X�:�椵u&�w�.rmi�3@Q���3���d� Sġ�!����in��� }���L�&���-��a���:3�"�2��F~GcЌ���|�,�Հw��,���c��$�bz�
�N]+��8ݫ!��ʡ����{�yk4�]�RfGЫ�����:e6F2��Þ.DcS��
�&tO�b��*�!<S{�
-�+��輡�p=�~{_B�+��)�\��-�.J�����־�?'����,��p����(��9�̿9�,sU�t٢�4�;K��o�)׬�+���\�1��x�>��ʐp>A�6�/�҇y K������2&K[~b)����Ғ�at6O��˻Lih}�1������D{x[q6?6�G�-a�ƌ2ꘉv����p�5vl���uW(/�%������ϰ�i*�ՠ��g�fw��]�A��Y��\��=h4���%�u���1��&H_�,�?K����ݕ{Z���.���Mf=;3jX���������&,��e({���8��ӑy5��b'M��!�⁙6dգ�'R�����n3��������,[�����.'��\S��������z�k�� 6ch�ؐ�,��]�댘8{t���ȿ���ZZG�@S�j��ck�F�1���<"��-UY~7�농F%O�a�z(��<)�TR}���[���m�7(۫�".���@30lҌr$D�_��E1�4b6�"S��΀^[{��O��iU;��p$lkkʆ��d�["kX��q�#9�s�L��2\��v�
��ŀ�,oK �q�R$M�`e�u;��l�*�i�ٽ����ߵ�V�&��s$�Yn	)�7�0�9G��T�ڰ�3�����0*�v'T��|+�஠��Gٱɲ�ar8/^�P�!���k��5���*�8�� ���!b4��� �x��x7F�j�y�V7���o������aoJ��y|�� V��ח��(�0��N���x�= 8��F��ǜ�<Ĥ��S����O��3�#�Gj��;G?ߏ,@��y�Ά�����Lrqa�|���@ܲ�M)�=(N*oYf!��Ƿ�TL�r�d��6�k/���S�_4@���C[n�K*�ɍ<���]�4����bΖ���t��*uԷ� �G�'�0�0�ﰨ\?�-��³����$8@]jxi"΁��5��7[F�G�<Q��C�ϣ�X;;�,���.3�~������Cc����Ny��QC���U���+
[3;�C��S�ӂS�xx>M��ݲp��cW�f#�9��rK��G�Dp��d66��}�]M�<u�.�q��@G;^m��9�T��Oi����C*����y<�=A�R��V� �z3��_�.���oɋM���L~��`����\����
�u��������5c�g��=v�����PSDr.r���ɓnm�}@�}&;�#�����.
�sf���2��r���Y�.y$1u�D��f��z����0��r�y{4�B���6� z��~��)p
�JG��n*d��iY�N �&��U�� 9��3�Q�.;��Ʒ����& �������/��k���M�T��%�fNOK��'3��+��GA�I�hڛ?���wJ�S��ͮ6������:�*�aW�;�Y�7�1*�����J���-�]��B����$�XW%c����%b�u�wa/����-k�;����_�hױ8Am?�Cl�*��r�5����s��v,e�S7(5���=K걓$���u�թ����Ht��8��k�ZK�"��~�U2Df�~���Q)l+gM�X�(�����i���[7��c"լLЬ
��U5�wq��ۙ&JHӍ�çh���5���o�cm"��	��`F��X�k}�3�#\Uݨ�m�$jLzLSP�dՙNS����Ok��5^F;��}!7�!x�w�vSm�����z&Ȗх�٩rvss~]��H�$-bQ���4b6ϝ����V��(zϧŻE/�q:�Ə*�/5�d�\�709�r6T��,ǲErDt�OczSS��>�/����oY�xE�̾E]�80!2�7Mj �����p��(- 5ԁ{���"��>I�ĉ�ysb�/hւi1$��	H��3*��H%⛩=�՟��[0��Y�Z��zQ���0n�`<�϶�E���M��U�X�5���`�W��ʚi���N|T�J���H�+�$I�(�y�,Q�E[?\������|rz�i��!�3拚��Du�����I�z3��o��#-]OfafF�L�ʁ��z�9���e�{#�pZ�E��ِ�03�"��e�]��藕?�U�B��ĠU�Br�m�h��?bz	�����*j����*g�2�ð ��3��V����7��4-r�p}��Xi�J�	�IU�o%����uCc�m�MK��`�7�̟���L�(���c��$@5�J� ���H4`*O%_���b:�
`�ߛ�u�ݛ��͟lz���l���mȻ"^����C7`���v�����6�[�g�hg@%�Q����*%;[Ɖ�U�C���g�1e���2�����Q`Y�٦9iMb}��Ź��L¤��^8�H!��	9C�-�e�9-I�/��Q4��ژ7P��x�%�"o�{"��IkQ�VvMu�\T4�- Ԡ��F�M��ȵ|ev2�� �Ip�|LS���g�'�f��Չo�8��FL�GԌ��|,�ը�f?���׉��Pl��ҏ�?��A��_p�P��1��ы$��5,�| �`M��!�7�1n6�I\���b'q$��@d��DI�z=��,o0�ɭl��C�LT�R���:��o��vO��/�8C��[_�Ro�W�g)hhc�WY��l���ul;?���G��*�y��wo!`6���S�UMu;h���~rwV��\��Q&��	�����;��_�z�BE�H������]�b��(��]S4�66j%� �`��"?$� ֿ�+���D�szⲤ��al*~���{���o�>+�U���}��Z�!��9	&ᚭ;�4���Iꍥ3�o#����8R�ŭ:_�Ɔ��g�qV�>� �[DTcŹ�,&���^M���cز�
���=��T�u��\���b�"z�F޻j�k�n��1�0}��se�2{.�0�$�V�8;��)t���$��<�|��L�u��� �ѳf��@��_�����g�I��T#�d ��<�	E��0A��%=W�eIp�=-��Py��	��i��5�B��X����C��E��RӡF�@�pt����l��q�6�T��v��&:��e��|���':B��^�4oB��3s�FIT�F��L�=4$.DU� J�{��j�V�\^��������1+i�,�~�>���7��L������A=ñ~��C��� �j�تB�X	�����H�-`ަp�X$D���L��i||��?��蜮Jj>M�u�:�K[y����Z� ^�*}{�2p�S�N��R �A�� �p�i�q�n�	��2�W�G5�9<�!�^��@�?K����:�u�o1ə����Z�R���2UB
��g�:���R���*���- �.0�LDD��2�e��.)���B����T獡+㜟ԕX�?��دa@H&T�IaG|�[�+�pTe�R��|����#���/�^N��"�ҕ����ͱ�F��<m��m�e{%u���o�4��?vS��Ta��+�a��j	/�s�~,�0Ŕ θ��B����K��=��´�{.��J>��Xb�|�B	�����7,.MDΆ�i��qK�g0������c�E��V�c\;��p�I�H�B߆�����ߞGj.�%�à���xy l�)_9:�nc'T]��_0�j��#�=��K_%~=���Fg�њZk6�1�7+C.j4E3�|u8�g��6��	(�1�Ed��sM��|!�z3��`�y���q����������رX����6��Θ�Ǭ��������f�����P%��lVq��z����Sʘ˪$u��߯^�3�C��W�$�#yw�������vA�{�r9��F��8.r�����H��&�c)��L��|��خG�q�򚚢�ibQ��p7ɣ�[�ّ���<OFsb*V�?�y�2RG��@�76nOdj�𑎕� -q�>��C���o���B�D�e�v!j�H����A���q)�`���<��(�R�!�H;l�7G3H` gh)����Õ5�����h�6�p�!tO,5�-쎓R�=���U8��d��N�:���$@?�~7�����S��<�jM��|�6�A;�ig�I�l����"�Zx���ـ���Ҍ��\Cx������2dg��8�U ��Ї;��+����e���坶�wx+iu�oSZ�������1�$ɽX2\��[t�)E����{��
�);�;�z0����5����h4&d�*�;pR��Xu�O>��A��d��� ��}��F=u] L��\"�MN��3�TZ��������� �j��>�f@%��Q�/nɞ}$m~A��C¨� Ut���$`�F�E�Xv��qJJ8�材� ��Ǒ�8�
g���Z��h��PY�� �lO��f`Ui�,OmtU�4��H��h�<Av�$�J�'���}�\��Ӆ�'�����Q��Y�=щ��o�>���x�fH"4i�N?Ç�4�!lg�_��� 5�|bP�C�7zSvg���O-���H�f�T��噱���y�&���"�����z��( ��9�Q�'�9�p*���������_��&?á�'�T�k�J7A�����.0�i�Nj�[��V:`��E���gR�X6S�t��
�,������<;$����"�͛�^��O��l�� ���,Mmr.#��Ä-��bp�੨"�G�q���,孶��('�f���fu&����P]��|(ȸ�p��
VQ~��҅���eg���ˍ̹{�!R#��Εm֮W��H��t���w�8-U89�s�/n������Ö!�z�џ3�:4����B��"	G ��f�s'~}�ZLF���-G%!|I	&�@L����VϹI��wr$Mˌڢ��:�w:�_�g�� E�����]��h��[9-��������2���?�-�*6�]D���`z�e������x���Cf��<A;A�۱�ilO���S���g4��OmǎjŎ�h>�ԨF��?!�8��6��OX�&Ols��/�cv�XZXQK|?�VO�����;f�Yv�W��Φǂ�!V �5JA`[�؈��ޘ�5�E���[$S��HX�#�>
Η��9�?�+��즸���efr�:�y��u@	g��g����(�z	�kW�;�r�q��l+�G>O�o�ɞ��O�s20�_ه�t����L:�f�/�|�h��yP���pzm�����`��[��6<�?y�i�l�y�<���M�mR�*24��z yw���t$� �#)��mF�g�dMA�!m���Γ;$���
ۊ��$����}Q�K��M����#��:@uq���b۬�5n`|�Y�#@���������T]��G�D�l����:,J[q�l���D�{�6�۳;.�f�9��8~�D�u+��Zٮw�L�으���ͻ������X�L�҈0��'J'�Ů5�h����=Ie+��� �>�8�[�$��=iE9`U~�γ�-Ĵ��b3�@ܳ���ߜS�?��s<4�2"ucbS�AOb��#�����^ e�+il�uH��b��t�|PH�Q���퓚�;S�Q0�MH3�l�O�	�*9�d�-�	�"���J�~�ѓ���t{]���QSp�~A��T�+���✸㠿����o����}����'��Ѣ| 	�I/��8���(��vz1g_�&���|x�Y��ON�f6��u$�^g9-M�X8?�^1�</��/�_H��Rp<���3��H'�}�TCx8(�Ӧ��:��tgo��5N���y��՟���>�~���AV]�1��h�i��0�� �����<	��ax_�Q�G��s`�D-�4�d��
�ւP�v�y.�A
4�#D!zUv��^H&�.4�����|`M|��*�ƫ��N��0%O�� v�w:��+�W@ -]�r��-,9]���.�k�`W(Q�����r�z�ZH�	�6�r�1��$��2��su��Σ��;�c.�G���c��X1>��OT��8'#�\�Jg��=F�'������I�la�}��6P ��w�[8���3�Ȭ��&%J�������(�l_�rZ#�R^�S�{�J����̉Nb���q�ٲ7
2齷���]����*�)_<c����uS�r�yEV�@#ͮ�v����lh�׫Y�'p�z�̃G,��{�C�S�LhF%���m��ȒU�
��Y�R�>����^��@Z��?�!>w�L�M��υ�ݦ���n+���Ir�z�s�	�����G�T�J9	om���m������͟B�2�ẖQ��o";������v\����DP~���(��!(֯l���B�#�	c�x�����6�_fD�_��~�!��
���%��y�W[�8"pbo��hԿ5j��tߙ� ��Y(X׋V���%���b@.�I���^(*�Eu�m3_�^�`*M�-%_PL�ɫ8؉�|܌`qw��y�(T{����b�@�M��SǗͻ��؉����V��O����8�a��c�K�2c�ۘ|ɞY!��I� 7V���q�Y���v���'ay9�=�ruC����C��LL4P}���ؖ��� ����P�'As<9>cח�PW���
��`e�A�=����{��\��?���/fG2�}RBT���{$��yl`	��=�C2�����>�K��ti�d�sFy�^����|5�w�/@�,��p(}�|����-��7���������l!Tr�9�u�9�PU�1Q;�tx��P5VM�B4M�1���;+�mg�V#6�	h�
�ߩWπɊ�:�O��	s+2����{8�0�G�iS�<�󢜋\�m��3{[~��2��F��t�|��,�b�d���JW�����P��� 8���}�����;J�b_��bM��*���uː��7�-d��@^���vZ�D�-���NX������Pg͖����&�
I�U���YY)�R��5�m(�հ*l����� F.W�H~��#V�г� �uZҼW�����k���(�<�������ܜ�]�+ڧ*ƀ�S�'��z ���gs���e�3(T��M��\�9�߱w�eo�\��,��V��)�\��������24m�Y"�������ɺU���7� ��
%�`�8�\�7N[���DA%���iG�F���u]���������j�f�3N_<�C��`-����^0�Iv�e$�6~ӑ�7��W�B4Q���g7��7ik�4���~f�=n�r�x�f�&`��;	��l���1�1��b�+��QU %�zY�"?�2-{1��-���CS@��w�!�,n�b� ��|'�:�j�,����`�gIϵ
��~�6S��7���P~8�-!�=���֪�BP����
1��m��U�l��(g76'/�Ǐ+���Z�nd��r2�òe�v�^��J
A��4�!b���~��.ڴ�j"�������(�Ъ)(�:��U��F<q�Hz��Bzu7� ^�9Ӿo��:tq�~	�CI��#}����s�P���f
�q��X'��,=JP:/�l��$�Cu1¶g��1!ڐ�vz�m8�OHs=��g$�7PO���1&O]�V�:˗�q���O�W�9�R���X��J$�B�l�T%�NU��?�uO���AG՘��/0ٕ��=p��y�l�s��n=g��v����]|�oUIߖ�I��>p&����\��%��`]�V��v�'��ƴ�uF���i��aܾ๐s�:�� ���\ ���v&�S:�ua�d�7J�H+,���ly�T�?�7δTOy�F�p�
)? �ura�o/:�Ub��_9�yKv~�a��5+�Dݙ>�z�A�v�)�fj�����f���t�.���PT�IB�rbB��9�|�j��u�Qp?Ppٽ�_Qf��7[l!�4��"�}M��G�T��CL�|2�l�+��]��8Re��N�Ѩ,��`�BM0H�Bd,�)��Rţ��+7@E*Y�_�م�%�>��D�Đ�B8��L�ckpb�삯�%���W2�M��@�ѹ���x�^��V�{�T�Cs��;�_C�5==;��,��/��}*)�'�_�0H�D��v_Wrd[T�1+��c�������;��!�Y�ޔ����ΐ�(��fJ���MݎlUY���Β�S���E5h��������8�1������#��'>ĬA'�Bǜ,�GO�S��r1^8��_P��h�0��#�l��:��c�'��Luw�Mv���/є�<~���ήX�d*�넨��yw���?��LK��Ɠ��~���=�O8=�n���^L�1�K��$4�����L�7�gTw�8���`�?�/���������a����ALX3VG��Vu�8|Q���b?>VeqJEE�����V@;�x��Ғ��z��X��
�3v����u"����c�-�pۮ~|�i�����@_�s0֧4������l;����󁡙 �=v�����	������nTGA��w�!ES�����d.U�!��7l~).�0���K+�447���͒�ES��D1�!�T���_���~/��E��"��h���itX���k(V(2LQd��M~<*b�O�}ࢫ�]�*�a�'Ğ��7a�P�K�QδX5!���,n�;Xh�+�y$��>���c�lr=�Y#�݇J�E���)�+%@s�6��)���⅍�{��cb{�Y�� 5�`/����>9��m%_�Cs����:�M��YΧ��[%f"��t��6�[�X3��)����O���/.��p��8�^�E����r�eK_��X�
��R;%�VW�X+Q��oț%{�9�J]JA���j��Yx��1&)�PB�V�ss�sѡ���Q\G�U�_�*����l�{֞t�M�ԕiU�Y�RT?9��bg6�i��I���+�C��:d��4l�~3�����2lB	��if�f���]�;0�G�(yU�b+�S2M
�R�M�Aʵ���T�f���FC���V؄��ڕM�W�^�m���.�IM�U�&�C�6��D4ZRv�8/!p߲8���7����|��^��=�+tO� �$ 	奧}A�8ֱj��v/K�n���(��d�C�䰿T��������Rʪ�߲zm�/�΢�dm����b�Y�4o�IjZ�N���5���ú�?�h���%�?e�@QB���\ؾa����dˡ��k
y�R����pQ��1��%]����P�d�('!�(��!�rro��rۓ~�D
Z�61����e��P��Ɵ���s��]�1�;z>IH`�N��2�$���%�4����/5>�A"%���צ��r)�W? =n�/k���/�C��>�*:h`�����}�UMq��>��]����6U�!����]��]��@<	�d�v�-���S�|�z�g�څ����I>9K
s[nʒ��"� �d����{�;�8������4��_�����&-���	;���BU����Y+
*���-�B��e�{̱�hg���B�j�Q�W�<$��N���Cy� Z��x`c�Q��_�KY_:�����T�i&���yms9�!V�݉y͗�+&�����ױډ3���-GXj���N1�ʲ�)����/�a��J�~v�T��w����d���r1p�m�F��Hw����c��==��~%\���	 ƙz��^P��f��hJxO:*����Z[�1�J�w>e��%έ��~�,ɇ!�#i5������v��݊C��|����µ
���%\��<�ĉ�vl�H��j�3�A��MB�Q�u�b8���M,�y��l�L�����_9��E��O���ǎT<y��&�|Q
�d��(�%T�R��a�؇���%*|+���QwPI��d_%�_�ȕl����h���`
���h�Q�	=�@h,-���z��S�fώ�0��N�?�nÚ([Xw��J�,W���~�m�|��n�(��M�� �z�CԭO���;#Nx�Ҏ�#��U�Zi�d3�!r'~.閧��J������γo5�"�Z V�Ѹ4��Br����]q���`�
W�-OPmƌ�0]��`�8�q��O�%Y�6O���W��;�v藤�Qo�n��;E
����&}�~o#�N8]�h��!���n���O�ʡ��/�,"K�6���Pa�!5���(_�9�{�8���i
#�˒jr�����.��K�&� ~X:�up��ra���9Fv�������j������l�e�65*5:�_m��ak��R��fs2�3N�V,{DvL]��O���Bq�M�����6�`�qűk<�\*N?�������A=���!������yD<[���g���h�T�藪u#�Տ��Q�F��z*2��z5+�T=�7U��U�e,?��nti��Y�p�R��kV,;�ER�"[�'����������r"��r��K��?���m�߃���p��H���'���@ǒ;����#;��:1#��O<k'�5]����u��.�nr�q�O�
�t1poג说u)E���dVHq�[ާ:< �g��6�s8Ss�2�xFp�L8�<��Zt9���hV�r����A��s �����S*ܞ���u9d}��r
����Y��yˍ�B^9��Ά���ɒ���6]}����nò�ln~����~�5�k���Ȓ���l�ڒ�{��Ǚ%soI��^��P�U�n��;4���a�U���'��h̩++�C�N+?|�<�l]hG�&�����Ɂ�k�p�!|�<�V|�]��A1m|��쒡;�@P�����Y�͑4���8s�K�%{;���4���R=���	�L|��z�p<Mu�y�gj��(iw"DgK���|�>��6���+T��e�Э)�u=���ҩ�&l� ��ip��~AP#�! ������9�E�.x��S�vՈn�"|S�Y&�����'3)��')��ц�bi��,ɋB�PZ����e���Mn��(�7H��t`��u��As�C[��D�D��^>��JD�A�͜�qE�W��Cm��&tL�$��I�A�����������4�+)퍿��V'�V�\�.է��A��K��Z�p�.Pe�*�^�xL� ��$�n�'������fZ�. ��I�O �Y^����ie���=\��^n&�=�5B1ĵ;�;~���s:ʇ�nq�9��ｬ���e��*-�T@�0��ǣ�����y�/Ϭ����iK�}� ů5��B�t�&ў
!�9�t<½���O$�������O&I�ETT�	��q֠��\�îW��YO|:2��"c���Y��
�7ޣ)p�c{��ة4s�Mx�e���_�9�M�%ڒ�\/H3?�-�T���U���2�������-���/�,�I�&�NZ���hQp�V����2��Gʗ^�>5��=o��dOtz��C*yį���Y�o�\�}��T8� ��`��l La/{e_�?��t͒D6��s���_+D��L-.�t�O�	�G�1�g�ߥ��վ��\�����᎘l�'�� C���w9��_����G�\�}`���@�Ь��U�Mw�����ʧ��J'xS�����Iyޔo��H�eҟ�'��`�9*���Y8�)B�Mh'!�W��
##1�W�G�$�q�����ʐ��~��`��\�]QX[ ����X�$�Q