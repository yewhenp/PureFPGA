��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ��%�͉�ao��u��� �z��8�Q�f��_=W�� 
�l�!�i�n���MK�Y��!u�<d^�2���$�Sb���/?��;\,����5ܲ����z6�����%ۈ}�?��eu<m��P�ыo~����z3N|�I�;z0h�+����m,�/�C��Ҳ�7s}x�p��?+���W'�@!Ɖjp
qq���:K�`E~Q�lG�`�g�H	ݒAȡ����	~�}�337�������G���s�����eۋ�,>tA ��u�֏����⟷�{��Mw���m�T�t:���3���r ��cp�ĵ`-�B�\�K:!�ik?�<]b��93��[�'Z�C(*��+ ��O��ڏ<n	쐤������E���l�E�w)��Zp$R�5A�FA�h�~���6J�J�_�{+��̇�0R�U�k�U�6+6�)_,��I��������)E�+n���`HeZ��<a���RUu�H*{�9����ĕ�hi��\��K�n ����h5���*�%��A���U�ԁ�#�rܷ�]6�i^_Fc���L��~����Y�r�C��q�k�wji�tcɟ�.Ǣ�b�t�Y��c�)HEЄ�U�hs�9�T7Xb�S�1K��x.h"��n�@�$1�<X�@�_�T΅y��[#�.�rk+>�x�{�Rw�E�a!1�20eT�LiL:�r<6��B�G��������
�j61}.�F�|��);O����Mޫt5���������-ؕ*1x�����C�����P�Æ���/�t�L�F�ae ����<[���9�ϞV��}�GQ���<�L��76:,�>-c��v��6�v�́� +��&!��ՙ�jsZ���`"�M:~�~�NO;^+���ⰻ����J�,?�������%�|��~��J
Ǖ�Tekqm�O�v��ZW��m>,dt��R`W*]�̀�c��ΊE	�U�Rv���ﱥ��<��"�W��#N��A-j�W���>����GI��^��( �<�0ĩ�%a1�Y]�Ь�j�~p���C�&���a�����?(�"E�۞Ӈ���m���s������� Ƹ��-�x�g��}Iek�&jm�� P�[|i�k|�Q��~�L�B, b�hQ���.H�Fʨ�L.��C�Z��Jܨb���O��h7F�F�h��.�I�X{���o��.ºr5��)�)2נ�B����{.�Q�}�e/�����(�c,P`l*���6���fb㰟�XkӖ�����s�Ҏ��Z�쵤�ZYzԃmb+�&"C1U��!����2)��g�֠�5)rE_ӡ;`�-�R{�,T�������wz��%e'RUW���:W"	�{`/P��h���򷙭���Q�n|�B��:�Q'�F+2�����`z�v�eJ�(�K��-<��X�8n���c��yL�7����#�
��N��Q��|��ٛK��n�(�K���&i����ԟm��$��H���Y���zќne�����F�X)V������/�Q�3/�	�ƻ׳8x5���TƸ��|vF!;唬�)�L2Q�	�!�ba�h&O���b7�`�j!5����s,�r"� .�9�D��:Q�3�w�0��m��mpiCB�o)���9R�l.U�'q�u�����}����aqz�9V�S� �]n��pu{���_F�,�� �R�>���Rl�]s�����R�by���i�10��+�J-p��a�X����kۺ�����G�w�=DG2כ�������V�z�h�ƨ����k�Ln���OER=���I�9U�� K� ������X�3�G����3eR�Î��Vj+k����{�J�vi*e�\j�}%��)�{���=-���jA'x�c����+ٔ��底rk�:8o纍�5ڲ���٩"�:���x+5�_y�(z��RX6���3F�p:0 v�Q�B��`�{9�wJ��u���`0)�k��IN���)��3�ն�l��j�g���T���乬[����jO�2U�:��c!���0���=sZAY$�A���5k�!
�k��G��g�E��w�L[Cq�pJ�lu}��F)�]�L�����:V��Ęp8ᩇ���1�z�wrɯ;�Q�G��v��-	8/��A�L���B%��%�+M�9�Ň�s��em�D���=<� �F�G�
1&ѣ�5p��~Ϗ�dª5��"�Z�F4�87BZ��uh
%�$�������DÞ�������.��LVPu������'\�A�h�;����:,���?�g4Z�!��l��<�2ܟ�,�l�3�f����f`�֋FW��W���HpV��9��>�U���<}�,$�[{S6Ç�Uvـ���V�(^�G&�B1*���0Ne���M��B�I:�3�@,_.
�	���p56ս�xW�W��O�P���X�_&��)���0��x���I��o#�I�6��O[�~�|�!��A�գ�1/%����ڷ5���0Q?gx�7�֕������O��'T5q�o���<H����^D�~�(jY?<?���Q����?q}l��{D"���Ӂݸ��;e�VVm�� wؗ�s{R%A�a,�yAI��݂Ԝ������?�a���$�[z=��c&z3IP��K>)��k?�9�/w�~$��z��գL
;�yϴ���DU"3 ^���<W♣����1Ӥ+Fne_VāD�z�t Ǔ��C�Ǐu���{����1&9w{�����xm�M�,p|-Ьߥ��yϩ�N����~�Q�g�C�������`{�v�h�l���`�m��ᩱ�}�R=|��!B�R�w�^�8@$N���?j��!���#2���ȕC�4>��1�z0=<�[T�����]8��у��)�[��$��ŝ��au9��@�ödՇ-9���;͍5]�Bf;n\��(]�Ў�[�U�-�4T����g����L�)2)����vSɴ�GF�g�t_ ���CZ��k�7O����n�3'�{6���W��۞Gaʏ.��g+a�����>U���Y��>I����`��b���a�&;T���`�qnA5���^�5^'��IrD�Y�m�{�(k���"h=e9���� 픊͓gG��EFJ�m���������e4@?�]jc�����}�	��D^d�r�2�wD�(�O�� ?��%:C�`�!�Ԉ,/l&�ŋ���A��Z���,���]��I�H�,�>��A��э���Ī�u��..*��h�7��E�9���!�U����D�����q����~�)~ܢ�ڨ��� `_�g��x��O��;T��Rͽ�{��.�f�(�_R�wr�4^j$�;�k�%��*��뮫��x��D��)p� ��,5pz]�<3+���#e��%��A�B$�ՙ*{��]��Њ4�W�iSW��m͝l][F�����������шk}���p-������Qj�;���b��5c�A� a��q��f�k��6m4�����
��K���j�_D(H��yA����X;�0\Nb�<�+�U��ݚ�&�����7��52�F�m(���A���:=ٵk�{D��N� ��K^i/������Xh�n��h@v�7(
F;s�کa0q��_�Z!1S�Q��J�o,�J���#�2��Sŀ����.�Y�Ϯ�'�~����
(}��X7�8hK�;^����R��%>��L��Ќ9-�i�&V�~����t��@�XӰ��4��z�mv�x ����PD�|> ��5���=�"�[�jF_��U� �Э�>�f�y�^�`G0k�z-�Λ�s�H�J!����ȌH�M}z��d�(_Ym���{s��}� ���ԏ�o�9�(���+��\����Age�MyR���������j����2��X;C7g�R�'�����.\x(��.�S1�c"�6ٲ�3D�#���B>�}=$�j�d�,OvGÄ5�hy��\w�F3��Ã�I�}�QJV���C���mS:��H��HLNcm�5 �D|���#��"twP���3���l��{A�+B��S�н��ߓE�Z�/+<h�9.i�3(�Eg�װ)N�A���.����Y��&��v��m�ǚo�d���b��4i���eĤ�D�W���E�"Q�
K��>��gQ��a��x�sI����R!t�&jG<MgJg�g^Gj��3�� T�{�$L���R��y�7�e��Z�����kI)��A�e��_t���`��(4����EV
�g�j?2Qz�q�'���' .uj�*%�k��k�)Og�~�#6|�L���<=�o�[N����s�bB���T%�s�U����7;F�3Iܜ�T7`}��L���a[�A��X�x<���㑣Wz��Ǹ�i+�o�E��EL�G,�w'�uf���ǵ$��� VՒ��hM�6�P(�h��@�Y���D�ε���}��[웫�&͍�{�5T�u#�Ϛ�B{M<�r�

6�\��L��e(L)�v�c6�� �ZU�.�,'V;Y|��m{l>��+}��#�����h6 d�}� ��?&.�۽�؟��lS���e��8�ūW�m?�xN����`�
�|Y&�j��v+���M�7;��ۄFeJ�����#8��qp�L�~僡���OC߁�"�N�'{��KQ/q(G=)y�-h�{K"��V��S�w�e���8*�����q��#٠4��p���L4�\f7>8ed���}�A���P���x�M��	�~��f-��2�����\��B��k�u��pX���:~�Yߧ�nBL"1 ��ե�����h��+-�oZ�Z/PS�dyǽ:>P\mdEt_`g�e<�^�t?�[���x� R�h�fa���=��-"�ռ0\��|��D`��mm�CİY�Ɩ�k-Xq>�dM�E����ia�;��_��ck��W�%{�pM��S�'�`��q�ۃ �������8�±���Sх?�n�F&�n@�β��ew�6l2�ɳ� {�0�(��^f�NӲg�D�k�|]�b��͉���P�y��w���Y
=�d�Г���sr�L�I��]��Ӆ��Q@��U�����,{�rs3�����ը������f�.XhIX:�)8%�i����i~UjL���rY�zZ��M&�F�~.�5�Z*Kfx��$�>������!#9W�aT�<t)?�g�A�Iw���=����oU�m�@�
Y,�a^��h��m��J{��ޭȿ �v�KW�^��-��'%x�rG3��eA
y۳0��	$u�iX��?�Q��Cw\�4��~�i4.m~�<��gT��[G#��r"�Z%���AY�f1����"��A.�^�>�crL�]��֥!q��y�]�� ��x���u�">|��PW�)|��}d2����x%K@�U�g��/��rҬ�'�ǔd�
J[����o\T��B�����jQ���dVx7plȂ��"��e������M_p��c�3��E���e�|P�������ŗ��E٧������ߏ�O� [�Y��n�b�򂭃S��PJF}����J�?p��8�<��B�������l!��l5�'�Z�py>�*Q��ׅ�>�f:D�����5�s T=��y�>��$�U!���2?>�j�˳}l�����+�����j -}���<{�,d�l�����������>���^Qg6�9<��Z^L��>���ߧ��Hǧ���F�����h���`�'#q�[C�*Xw�Ji�F�����DOH¢�"������~�Xd�h�����" �=[��L�D�F��b/l��UEغ�U����n�)��抇��Ь�|δۃ��x����{������w�[�L���WM��f�p�C}C@�P�r����ҋ28��#N��H����V�Z�	�s��ә*/pon�Qۓ�X.�O��(XT�R��z��7�L��,d��e��r�#3� vY~���*�N����J!�g�:*h�axp?�/@�\�ԃ�ʢ+�R�uj�W�g����L�,����

�qԹ`��	����,�je�P�p�#��h����t��@�=NR���W���Ԇ��ݥ& ��3�5�Â��;�x�g �:�ڄ��q�.�U��VLM˚�`��D5�y���_�K젫AAp1���_[�z=#E��H��?���6�B��Q��:ˢ��-���?c���������b?[��(0c�U�P��M����	M��:�jb"ߜ#���kncj+�SX�#�Ȉ���&Z�.߀�[G@�(���5r1ɼ�"�+͢^��7�L�nO��9E��I�d܌ta�'��"��C��p
��|M��@S���� �_!R���g�J�$�}UM��ȴ��L��ȉ1� �ר2��WR>G�����^�dx������"��?�n�.�l�xDI����C�q�-��1�n��O��@�j��B3ݙ�
%S<����>���Pb��c�� �6Q���M���*�?��fQW��(\�a��0��J�����-.X��|�4�%�Y��R5f4��II�&��TR��\������"Feb�i&��P;�ƕ�^� ��������%�S��ׄ2��;A]H��l�}oC��D}�C�.Ey�{�8d��֎�"��*6��$:�]9�!��(�e�AYؓ\e�����Sؑ��߅n�ˏ|�K���������Y���]����\LRe��2��u�|��Oz�����'��4^��#��=�QY�9ڠ���	'^?��ZRt ��K-�ǩ���Y�w��� &�������&r��%�G��w�E�����!�Q@������aHme�k��`�>���j���b�Y!N՗��ӝ�PPC=����_$���`{�ih��#�ೂ}�9�_S10N�8-�6��o&�
����b��9<��/~��ZS]k�m�IpGʱ��`�-;^�1�ͽ�@yb�:_12�8��i��T�����r�9ݕj�Ǽ�9z6�;���'y��-c3<�r q��K�wn~�t�����Afa����^�ExJ����-��4��QP���6r����~�S��W@#d�#�-��8{���+eRi�m��F�"��d��KIv7�A���5SeAf`�_���C�:�M����!����Y��Gfw�F`�
�@�E��x�����1*Zx��f��ۜۣd����?XS���iu��V[m�T�f� �R�s؊ӗ+\�E�̒��A�t5��U��Rx"{Ę���.�}���kM�o��Wȃ�ුM�:Z|�� A�h����%-\%(��;������}�6���)��;�\]Չ)�5ݢ�Δ�b�ߞ���'��:��ކ������� 9��{���'�>ˉ����ݱ�?[]U_�����d;�?Ow��W��O5���\�TE-������e�[M��,G�#H�W�q���`����!���5<'�b��]�/<�ʎ�@m�W8r�l-1�A�d|���_ �O�ƤD�	�r�2�a�1�>� 5 w��ck���_h��@u)��J��@��3��꜔N��u��}�����)���K�9[ƌ�bcC�^cc�t\��B�P��S2R��β���:�*�,����(�e�<�n�^$��y��Щ��a84�?���8
�	�u��1���Qد�:���������i�a�p����m6�^Ҙ��x��y����W�����������X���ݒ�9g\&&�j�!�рȣW�}^�]O�ِ2Ɲ��l����ZE�z�Er��Xy�,�*GP��=.�mz[�/�]\�ȉ��i�B�hs4	����U/6�T��?�φ�J��C�(��'~W)�۝"!���ɳ_����t���ޑ�T��ֳ;�������l�h'��\XG?�ב�`T�����3F'D������]��^�L����^ ����B��Qf�s�#�&�"��� l�4�ǉ`nOdr	��~��A%�v<��K��1���y��)�Ḳи���I�}z����������@!��P�1��/��M��9�J Z�������Q�8��ˡ���T���&���qpImI�wJx{���z�0��3RL��Of��h��1d��盟�5r�K���f�As �O��K��>� ���,?xSR�mcG<��	�G��0HyJ�����B(����#�����ጩ��# �	Ӭ�(H�vQ��83�gI0�4>ب�r^�$4_%�;st�����o��tz�ؔuu��!g( :,�P������ ��ue�V�����ԩ ו��h��.ejF޸s���$"3XM}���F�~�1=?-WD����VÈOsl�2ƀ�� 	Vxv�>��
L6����,�	c�u���9�'G[i���D�����Τ䵭��$������tQgu@ ԣ�=a��6~��1��_(�+T�J�ʔ���~����Ρ�)��C�@D44lR�\��z��U>��&�S#>MrA.;s�6���fM{w�j� /�~>�I��;�}#�Mhٰ@� �Sk��u�oh����ܾ�{r����"mP��Rd}J��c��Tq��f"T��B8�����nNc�?�)�V��/��0Sߊ��=� �D�1��\P���wx_������{o�Oi��~�{�0��Va%h%�K	 �Cæ����}v�E1���j���XM�eڀ�t�)���+c����^^G�ӄ��Zy'��ƪ9QZ������oEN�f�h;�L�N���rU|����Gw�c�nɊ���v����|�tnf�Qz@��f�YW�k}ڧQ6���F���Ym�$�&�U���u�GQ�(�'��P6�+ڬ'�!j;�uf!����L�o�۳O����!��n���b%`:�X�Ed	��s 4�I9�⢮e�m�){XB����;p��4'Y�����.�D�vF�0 ��JHD٣�@^O�O�!�^�#J��iۓta2]�R¯��_ ��!��R��` JJ��Lq'<�+2��͸�_�p���64���'R�m��k���.u�B�)��u�G.J�� �z?����&����p9�x��ߦ'��V�35�DΌ�C����Wԛ��u`��Z�͛o[D�K�}����I�T�~M<��V���'��C��uU^�۝��J6�H�"Iז�u�?����ӫ>+_e����A����Q�8n�t�VS_W�xG!��2ewQm�-��qW$nUg2�$�e���E�a�<S����K����+�vr��b��(�X<
h_�c����У�ѡ7Гg���f��S���C�&���r���t߀��!$��$#/��*W�#�83*��9VTϸ�|�E��^��F�n��	ߋ�r�|�է�SPzG���TJ���)�)�����v���<I�,���C��U�+Y ���5+����D�\*�7P�W����\�$�Cٯ�tW뿞^���C6�*$�� �F���#'x�L�Z���g(��@�Ή���6�ɪ��~��Z��O�6�8�Sc'1Ne 6��d�� ҆��S��~�cn).�����������n�Ь��*�����'���͟�QK�Oǧ=sˋ�#�b��5�.�o��I~r���ME }zԼ<��� b�^E�t^Q�(��k9\�����} �n��?�����뎠l8V¸={����
�~jq�9�:�;xg��٣Q��{�P�hlɤ)�_uМ�OS�\�_A����@�^�}�>��v�Y»�x׹��0�'Ю.OxUq���d)'9 &s7����|���dV��ٖ��Q�u##�tZnQ��v�w.��O�����};�7�C�4}6!���
�d����OЏJ�o|A!L�޴���ȗ51��H���z�M�z%k�����E6�h
^x��B�E�f�P��J ��q���m�9�rG���gn�f8�#c7�BzzN��U��qS�8�=�ӊ��9T��E���;S�l�7�����HM�d�I'�4q�u$}8�h�
����=t�����x��wAey#�u�B	�jaR�����Y�������r�
���&�@�����#e�}v[8G����?Jc���8�Ǥ㥊�02Y�3:V�۔0�m�����S$R:U���N/	�ٞ._Π��?^���j;E�"脐z�[y�yvV�������� v��.� �����^'Aq	P�v�V�ㄝ��X�c7�S�H��w���u`A<_D�~˻W��pp�,�j}����V_�`�qi�]�8\!ܨ2��P��Y|M��`��߂Pެ���F����<s��b���jw�����!���6E]�4�'4��6{��;?�� F]����Q������8|�w^UW̻�x��vG�Ĉ�[)�����rW\�2�R����۩�K�n��Q�i�VE1E�谒oթ��'�)T3�`�E�_���S�b����~��ip���,]�:����j(�:y���\�
��`�"K�;/�Uk
���ZN�U�F��i��i�L�d�Eي1leZ\��pf�>��h�j�伞�7$���I��P8��j��B��6���?��W5+ҕ�	��h$c��b;���o�=R�6�~xV�L7g���R�&��gG��v�F�k$�v�Ӝ�B,�7�s�O�~o�)��c=l�;���e���{8�����ϯKb��e��0���� �,��SL-���yy��g�+��[��QN������%�_%��/�x�7R�+��ں�\5�ט���������\���]=e����RH��4]�9/�z
��K��r2�R��om]��}W)�m�"/F����S��aB�+�;JI�XQ�g��������Z��A���bx8U�	��^��q������rpO�ѵY�'��'���9�}:�~�"�
_۾U��x�~�ͫ0F��Y�A �V����vⳘ.���K�EvlCRv����ng��w�R��Δ�eɬ�hn�"=�]=U�-F���ψp[��FW�*�ac��_G���T���\�ճ�u��A���T����eL�� �x��L���� Fb4?�~*ڂ:q��nf��A���?s�7����0Ɩ��l�_%l	���փ�w��2L����дܷ$J��KD����;��1��r�7�������������dm�Sc�F�C�f���V|EE�F�����F���2gbB3P�`H,_J��H��}�쌟_<K���|g�h�TĨ�)f�t&���!(R�ϭ�J�)#�c����FOgx����
@۩���\���g@?����"Ȳ�J�){֮>Q�	 ����t�������]��C�z�GNc���|K<��B�?����^R��Q%�#L}�!�5�����������֜��-*}�0�0�)M<�>�Q��bs�L�[g�+ГĹ	,��2���%�jI���W��}��?�M ��j
��`��F�5'�?%r��6u!��c	�,��b��O#]&,Խ��7U����4@%��Wّ1 ��u�����֪�?�3W����p"�j<3�1�?;+� <,����Đ���Û�]��֎O���y�Ո9�V���Mv0r THz�X�^Z<f}�א�dȤ�.c1�U�]r}�@�
?.\i�c�d�^r���w�w%X����)�.Vޜf�����RJکA4��7��a��� �Q����|��8�%��D��g�([�,.�}��-�MU"�/��#�>��$��J؟L��<U�5R%=�w5����'u��BZ3_ݢ"G�e�\M�^�sS!�:Ǒ�I�����Z�� ��u�Q��`�8o@�)�"6*^J�B���^�V���Ћ8Xj �d�N�r)�V&����9.8gmU5�)v1�u��=�7�����������q��Ģ��c�w"�}�.��O��P؏�C����`ȒL��[��S ;?������N�=�KXmS�c(��{�?9wE��w�!O��l�l]GG&�]�e)�}���W?����N�l��,χ�Zm�c[{��a�s](:D�eJ|/[�z���=�Y\{ϐ�y�>�9�a��`%�~��2����텡�}Qmn��k*��ؒ �B�7�É5ȗ�3$��ځA�Id��n�!�R�oq9"�&u�E�X���9+D�I-��z�Ý+np�x����7����ȐFq��C�C�2� �Âj9;_��tZbw�̆���F�q���`_'��(��q~�����-(u�ob�����1��T�r���ȑ���Pp��RF�ߨb�og�6Z���' �þVo�S��J�(���)�A�����A�=ϰ1r�+���W	\�Z�M�a��[_��H��U{9��u���0ή����� �W�Y]��Ɩ�W�e��|	Ȩ��c��*�Dm��	Z�O2��o����F�j����0
Oܼ���'4�/���=���k(��C��nO0MǠ(���ۘ�[�<G��x������8�m��ܓ���s3�Uߠ(��#����^R�'�ʺ�q�L;x�J�����]H�����s�W�HABm8pg��P�ۄ&Aw����k�>,J�ɯ<���ᾼd���^��͉p�y,u#�b��vp�j�l���Z��R�lT� �����_�OK�]�́�(�}Їo��]���{T��C����k^��/��C�D�c�6�
,/4H z��ϴ���^3�PI�i�#��*��o}�����X?؉��褍9/ Z�Fk3R��c��:1耧2��*�q[�۝'��	U�g���z�����MxwWh9���W�4Sӥ��'fFY��N���В���ζc��t{c���/��/�}��^Y���Q`����8��-�m����t���т�d�cr�1c'W݆�m��E��j����
>'ϯ����	t���=!a���f)-�m�%BdWG7a"h��!�S���fU6��S
0�XH 6 ����E�,K���¥�H�V-�Tn2	:��MP�7�2��ER�1$���my��;��3+���y&���.`�Q� 1�*s�(�Ή��бR�輆�Z��8����%��l�#,�����sq>�DM5�{Mt�I(��k�8l�PS��m���_B6N�e&	!�.`�����q�;�b�cr���%��%�x["�eD���C;��2�vc�`�k668BB;���ȫ~ϧ��$+$�Ra5�Ī�?��vs��u9G�|�r��/�v�"FEW-;D�Z�~vK3��n�{��洒n����x�2�lE��G����5@�־0 {��n��P?�*>Q��u"����:�R��gn��3+��3����'�#�Ǫml��1^��\=��F&��4Yץ��PǱ�	5��#ƈt�ŵ������y�q�c��5��?Fd}����L۲G���m��;2P�(�q��;~�|6��$~�=7��ޗ���0����� I<l�q��?���[���EΦ���\��&��Xm��خ���	P����;�f:-�`7ݎ��I�h�֣%P�pzZ~�k�s��^���9�1mw�gK�
�[�@�][fD()�� %�aԢC�a  D�4��	M���
��װ��?���ʩ�ks�7�n#)��e�nS�����Eh;�":�
1��N�i]�I�N�����iJ�i3o}/��Y!��UR��7��b�[GP#�(W��P���(C׳��$g�xTD��;��$��e�C��\��i?��1r@?H��`�K���2Q�~��	9{�g��mB���O�����x��x�XY����0qS_�o�ܻ:���0�ڋߟqty2}E�!�;��Z�<���T�i��G$�Xje��ߛy9�ŀ�*�i���w�x?�a��N�d$�`�����I=q"U:�7�P`��E;tj�-�([�f��r��%[F@G5����^��)8oƲ�(=�	�l�[�\���1�jn�׏KӴA��x�)T�S��Q۰K��>}՗�D�����5��Ҹ�q�8
9t(ri*07֖SP>)��!O�n\a�aQ�u�`Z���*��X(�zq�_�?+�eG/n�(��G'v���	���C�m(+wZ�i��^�V)�Qn�yJPh2�3(B���ݎ��c�B�gQ6����io��6���8
F�"����ɳ��	J?�Di9�^L�3�K�Q��X}��R9Z�4ꑤ^�nRA=�Al��^�|�{�y����x!��:�_.��\.��6+�k���[O�|�qݏ�8�n�iV��_K�9�'#���9��X�0����f.U��?>�'��dV �!�S�bt���	�M����9�U�%�KMIk`��Ȫ+�Ԍ�%�s���=|�;(F���!��Ē9��`+tn����l�p�$��I#xa�?A��l_��:�"C:�t?��_*0��5���
K.|�w�`��\�F��>��z8�.��v��wU�ګ?�^�.�>y������<k4�E�"5m���;���8��_NwD�7,�6��(���w+��ܦК�*�,l+��WS�"��O��1uRB{�~$�6�VD�	([V�Z%��DP,&L#�\��b��Mb|���od��xN�T8����M���K��W�+�Ϫl���Y����2���Ә����']S��d9j2��6`*n5�>���Ҫ����`+���8By�q����`��I�i<=�UD��~�R�%^|v�F�'.x�����
��36�أ�՝��4���s@�]@[�VY�u��h,�t%�$moD���X8���:�5CoO�}���jX�9�9���A=�ɺ�R׾�ywaSʞ�r����)�d��̝��5�|w1��$�"���5>�
9�C�ZZ+HZ����~wX.�sJnP�Ɵ-��\'�2q����[�N��6��$��St����@�r���E� |����b�xӴ�D��[dL�ټ�C��L����&��7�B�7�s�0��rC��"�^gی��gJ�2�72; ����"$ h�ys%�_HG(&��p�y���ve��qD5�T��/���#�N����+.z�����y��U+�`OG{k7 h�9�=���%'UX���0��9���I_C�q�ϽB�N��D���mM��L�
,��2�Q�V�
������9O''�z�5��<����
l��R�c��n!�M��l�����ǩ({l�1g�TvO��q��D���%+�_�-�V�Y��1@O���h'5&��S*9n���eµ����>D�
��)@D��9����E��Y�B�"1R����'�����_
��ݱQ\��
��&k���� ~�B���5anK�u@ab�b��6�T9ڦ ���li��AH.�gP���kP��.�㻁7��3��pvG�S��]��h��F�B�E"x��Ng#�X6�ic$�h���S�?�E��i"���u���X� ��7b�o<�W� �q�=�&����"�q���ji�ئZ� ��,�{㧌� }W�N3ߤdYf
���|Y0ϴ�f�US����kR��ID�}L���í>n�aH��"Y[1f6��P�X�x��( q��uq}�R��H��d�<�ǳ���X�y�R΋�w��U�&�������8W�����(Q�xa���S���7��X�`�E?�A�)H�!%��ۤw"�3:����GV�Q|�;bS�Fر$��W<�7hB�(�� ?�X�X��*��5����8�\usM�P�a=�K�MH�t��ǌ�?�Z�<1�6�����?�s��w�[�����Q���:=i�
�.f�X��_�}bx�t��T���Փ��* B��S��{�GQ�{l��;�,�����_�뭃>@:a�w�h�;T������:~�ev���pf(�M�����3\�����d�ڂ*ۿ�l�����I�@Y�%]�p�+��U��sd��I��v^C���Ћ+�����4�ܬ���**��eA}èe�n2��~L�
37��ZNT�'�}x_�|�M�ְ���pi��"��	��]e>��q ��E�!�T�U=zT(���Vٰ����
�bH�6���p���ޱ���8+�7�_�k���ik�Ӿ�h�ұ��,@ڛ��v,���F��7� �*�`���S�@]�M�Qq~+c���j��"ίWTO0�Qp��_���߇U6(|,-:b���J��@��O�e�	3J��g�^ZM��:��l���t������0@&�B���z��L؃�����y��L��k���V_ů
b����~�m�����0d�p�=R蝑l�A[C�o�b&/9�;B��Ŋ��4_'�_}�����<�*����Zj�R��Z�MP~/����d��%7�kv��	^��j3���g��"�R6���B���+�n!�b���3��u\���H��o���3B�]$d1�
i��U�+�}��6�VL��Ͼ�^W������Rl���L�8�Z�D�����a�d�,_������~e�ڰ9�[[ʎh=\R�F����"���S�d�"w"]�*�l�1<�Z���B�x��GⶉB%��q,�{n�JHñ���Vt~r����?`���!��:��F��t� �Ozbǰ��oT�6O�݆U�?��txJc5ܷ��5�F�E}wy�T!��� ��Vs�6Q�I8�ɒx���z��Lڠ���wV+��$���cKH�M�Ι|˺|(Y��E�^3���(�dǫ�\�	aW
��"���j�����Ъ!6_��w���Ek@�����9	tU:ÎYI�v�Vt�W&�a�$��z�$��$d�@��j�\�0���vXB9��:�"
펰�3�`r�v�7����4� ��s`c��mK�!f�е���	yw0,p�hd�B�x�Dz�VY�i!)��0����\�s���q�y}�g �B8`�d0��W�䕕'�s��%��T$�7&��e}��P7�c��А��j���C����Bᔊ=YV��0�.N?0l��a(��pj1أ�Wd5������,zS0^ X��������/~�e�9lh����حT�-�	����AɁW5��@W���K�	U�)��
!�"�(Z�1��g�wT�*͞����c���{���5
ȇ�Ld�R�xp�>ˁ"Zb�L�L�.���� �(=�d��>��Ŝ��>/�\�$�]T5���	h?PTFp`�ݯ�ʷ�Dػ<l����u:f� T��>��|_���JUk�|��3�a��t�C�CZ+��ڕ,f��n?�m���ʝ}r��|�t7?Z�Op�xa�4y>O{_���V�3>�AL�6j����hf�H�����m�Y7k3EwT�:��0Oo�����T���NP~��ꆟ����&�|�ذ�"�\�΢o�s�Q̦�f3;.�0Bz��T�=����*l��7!�/�������*�}��B�S�xpk�����Wh��@���	6['���7�p��LZ��6���J�0��q��6B�k��El� r�?<ds.������q��I�n[��P؛IHc�~7(<��).b%�����_���
���->��gw��*��D1�v-70ej�N?a"�,ê��Pr�,����\������#�N��`������t�k?4؛�&mu�i���x�!��SN��0��Θ��V�����~����PP����VO}�������Z�p��y�CE����k8����|3�	�4Q�S�����2ơ�k�;]���C���H~jX���R5O!ci�a� ���[�|X��B�En����C��}��x�ȳ���:��@`!Y�6��CA�Z%?�>6 �ymo`�Й`�P�~�T��ކ�m/�.��%Cr(hM��I�]'�b ��CG�#g�4��w��F�)G>��.�}t�$턈a�/�F�C����B�£'������/z8�q~*��F�K4��Dnwo3�8���e�U��n�^&�'y��zY���y�^�q�b�p�9���.GG���{��֚¶�l��dD'��X�+i�l��ȋ����;�Ԑgz�Z8su����UW�Z����������A}�v���UKi��������K��%��L��DJ�8��32��>X�mJ��?��T�α�n�ըK�4��	������{D=x�(��^�"��+�m���y��:��_<�9��se���c}���t��{/\V�̪?�lG�eJ���haK���_m�4t��5��z�cw3�f��P��IOgL]��Zܐ��`������LxQ���^�P<as�!���t��I���j)Ǒ���6�����HA$v��`ЭA0���������_�׈�y��H!�U��K4kfٟ�e��2Ƚ�N��K帉�LW����*l�ٳ�q�!%�o (�ҶD��,#�K͋�ͦaM���+�ڥ�0�x�O�'��X����_p��j���Ҿ�!�w/<����͡�W�L��gsC�m�[!�9Ñ�<l�))
��4��=�ڃ�8�`.!Tm���%k���g�1�9��z�F������&Ֆi�
d�[cr@@��`�k����*Q�n�k�/d�Ur�Kztr��m�sm�z#�3��f��(�Qe�9%:��v;1���B9�J�@����	G&�4��ǁDP�T8Ɯ5�_^����2QkShg�nF� ���8T�,Xd�4w���C/��CA�VJ5�����{:߁�Me�ٙ�2@S��
鬗x�?{w���l!ج��!v�@�@�@�x/m��l42֞'��_�p����)]�)<�,XGv'�TBDT�x4"$+�����WD��8��r_B�8��mk������������a|���u������ݼ�������������	�9R�Ɲ=��V���>�W�G߲}WVý�>��YE����u ԋ�Se\�Մ$�I���D=��ׄ�t����_�V�J�*����Nʦ����}�������s[����k�W��t Fh��w�����Sp�#?�`FU6��z����2|���P1W�0�"	��_��PH�3��0W	'�8,����]+� H��2��H����	.���p��d��Z���~c���+r(v(6*�j֎�rǂ]�0��bd����\ �����Qҧ��OE�;c��[h�{k��}��KC�(�!z�⪶�*ohnCQC����=�zsO��bD����5�UH��X"Um�����9����\O��U�A3��&s�Eol5��y���8�q�ɶ2�M���\;���.r5V��U���[�F��+҃�5��wx�)}��d��u��TI�Fd���C3��)	^�G�뗈�r g�ΉE��L�z�$���?���3e�t��; $-�������|������2���.ʎ��_��.��A���/|%~:�l�ꃱh ;,��bG"�?�R-Ar�1�<��I�yI�b�y����6� ��N0�"ਣ!�s[���qS��8������d4�* �K�b�=Ne4�� +Gi�nJ��a'���+)V��k��������2�?�&Y,]2R�]i��ap��\F,C�s�����V��f��h"��������/��뿍���&�;A3_-������F�U��c�+�l-I�۱�oh����}C�j�V-+v��D��e][�
n	]�mK��u����/�<R���5t��u̜��G�&w�� W��<P���[���ApJ0>9�%����6���G��Ćî���+H�&�P�y��:��G���K�"�=#Pۙ��&� ����1��W�@� ^4A�l8Dze]�����JK��jĦ�j����!�����j�wᤈD;L���Ϯ�x=~��Ō��G����o[l�rL���c���ˍ��V���IaK��M�h���36��g��'!J�X������ǁj���e���\T-Զ��h��c��A�n��f�@E?�C^΢�Ǥj�F��N��{$_�E������@|���q�����ǯ�t��߂t�v$�B��(Ƥo�w4���zM��̟=p��"�o�`n��I�ˉn� )�4��o����1:�,����0�3}��/�*pT��߃1����μj�f#�_"V��QCr<3 k��C�e��U��x�I#����f�~���g�m�z&L�.xQ�n���!���w���+�C�E�.��{��J��u��<d�}X�ޮ*%&U�]�pڧ��'��|uI�8!t����V��+���E����4�RN��J
�-8c��?�e��Q��;���h���J���m�Dki��4��V-�/1�2ܮ1'dP�%��(�n|T��؈-�c�<�m�%Ur\d1&���Z�`sx(��>5j��tA�m�e�C���?H�ȡ�Mஈ!0��2x7Oka6� C�,wn�R�G(�|��12��.�����р��42r/='����>T�*���睗��"&y�;=9\(����m�ڙ�R�N�Hm��O���JSKd��u4,ү�U64@o��
�c�E�3~��m=8��ds�t�.�34��rh*o��g�V�F��W�aie���dB5��d���h,�a�Ҿ��n�9i�;ؖ�#�d鷿i����1��U��9Ya���K��׹Y�&��1��U���l7�ܰw��'�~�"�x6��g��sM"`<?�ŠLQ�z;:�
�b�����!�iIR.��������]�$c��k�u�ؠ�O2�7�=%�a�?6�m�����̔Oޜ��{�c�,�i�Z睇��1W˖e^�Tfd|	˸oV$�wڥ�L;ں55�(c��zZ�c6B�&.�>��(�
8����(bDd'e���k/��ȗi�����w����A���W�m����vH�� Ǟ�~��y�#���מNٛS��ca�3B��.9���y�]���Z"��;��p�xB���G]!����\4��8���m;!��d���nԨ���8J5`S}���}��#E��BdͩCm+�@cf)��WlTT��8��gK�Y�҄V'X��UB��i������|����3��X�!1[I�aA�xu0����]R��<����$d ˱��Xb0���#_4�Mz'uլ�Ņf��b=���I�e�u�'� ��B������C�Y����0J�I���γ��N�N�Cl��;@O�9�F��e�Ԉ�����Ts�N�Y�K{��*�B�}�zy8��HV��n�D?�U)��q&�n#�_ �e˜�c<�āxz�vo�,-ܿz�,Z�h�����R�e�g0�п�7w�J��/8*���k^�ır,S S�jL��R����1R����Y��y��A�fQ�&ON�j5�B%,��Ć^:�,I�XiY�<�a�馋�f�T�@��c�'�p@�\��mw�Ξ�3�� 2?t�����KҊYó�jJ!^���(�!�(�L0,�:�}8�թƌd����A��ROm_3�	c�����MO,����J�$}LmP�!o�V�G�+��jܫ�-�I�����f
Ig���q�X�y�Ȳ)�e��������8�D��@v@ܟ���|����m��&�q����~�r���}4�����X�0�������9���`b��%�iñ����]Pd����W�{��p}�q�)�іƵ��40 q�7A�Gr4EGiOQ������ß���~��Qj��=����i�V�ff�	2�o�8o��-DvǺ[�!N\�[����1��޾d��C��n�# b_u��;����I�dAS��D.��.���4�ꕼ���j���q�G9���w�N���jg�J��le����׉������ �:J2j$o�J<
�a;0 6%#G�y40Q&y$ ��E��6�o��($X��q�^�U��r��^�̈́ZT�7K�-��P�W\��o�+�#]	�9y�~��;��������y�f���I.�6	�h4ؤ_����D�.dKAt����I���Me�`�Ȥ!߿����S����`{�����#`e;.�Z[�f�cl���k��l��E�I�:������ T�X��&�>����Zk�T�o����?�Ij<=�ZQ��������=k�6E(��w
ig�����Î�M�v��?[��v�vܑ5n>��'7I�nh�ChŘ�_�!Ȧ����s�K�T/Vn��������_�������f~ە�Æ�D}�@F�o�Y�8|�{������ �$�ƁIxX!���P�l��_DJ^��?�������X�������/��:�}�.�v�ZW�f�@�!�i;�L[�Ƿ?nQ)��eŘVAւ3���ƻ��$��a��0,|���du��pn^���(!ĉ�ŋ����Gp_����hf�q4#^G�����̀(8d�RV��j����L42V�����RZ��y����_�4���jn� ��K��4�k�"�a�[lA
�x��ȳ�[jb�CԢ����YD�G[�����	z��xi�p�|���\�Y���p�O�\#9z<v�g��و�DmoW���C�X����ڸV��q%�O��r��b�|fx���(Q�����3[f�ϲ<����B�)ĸ&�s��k�)���=��|:�Q�e�T�.�ܑ��xK�j�"��M��6��E0�(Y2>�5v`�2�b��Z%f������Y;�p��l��<����e;��%諳Qߟ}#'(��љ~e�!����6�-�� �*d%=H:��}�#ns�<Owۊi�m�����!M��D̳
k�5����"<�xe"tjh�Ǉ�k���U��l��MQ�Z� �O�z ����3�����$��)�7�\
�@��/?����U�P�~��	PKYMh��p��&�X��.ʔ���fD��㮢����5r�#���X���}x�)E���T�dGί���\�k����pT��h����5�4N~�