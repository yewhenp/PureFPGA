��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_����]ׇ5�F$�,M�6��"�����hgu��:?)�V"*�T��2�6�v8,��Q�3"S�Ƀ���+3ӊ�ɽa�xw�W&���K(�j�G��O���9�f�L����?1}B_مV$�Ēߢ�3URj�����pX��I�"��%Մ@{���4(|I�`5��&NU���_/i�b�ݴ��-A��aZ0�p�,/�R�.��r�O���+��&����vqoUq�a_���{E��n���&+����'x��˚����+<t���zʨY�^9�p{DÈ!t0�-��Ò3P�gp^T&1>Qk�*����L,z;ғ�H��Yxz�Y���~�΁�&c��ȣ�g���*�l�B���R��c�!5��p��`�K6�jG�]�Q�_��$��r�e�T^$N��H�lN=n�-D���T�;T�Q��-���[��d��_"�)1LMʛn��|eͱ,�W������5���@N�C�X-��vz
F�q��X�(&2O�
�lW�c��r~��/]A�i�͎@�̐�:��y]mS�5WT%��L��Ыȵ#���ߎń�O�i���[�:Ix�1���Ho��<`u�T���g�i�D'`{�0U���ek�D���9$���-g������/ѷ��wM�6��R۞�YTT�����ʭ��&���� ٚQ'呴qI�����z���A�U �V�Sys(�u����j�%f�}_j�!9��������������6���_�l��\����T AҊUI�>�DX��G�t,�)&X�ʋ8�r�CN��A�>�)���j�-h��l�-�T��[B3�_qy�{�tlt����n����k6��}7A�PJ#RR���?(�I� �ޢ��v��UW���"��v2��2����2r����ku=�KnDC���M�rܔI�;Z����2+-�/ʐWG�m�*���IJ�u�ܹ )�Ӆ��v�����EH��Ĕd�3���8A&z�*�a�]�Im��	I��������/����ӌ���=/{l��:	i
�tg�Uʩ{�����q��>m5�#Κ�c��~��D3�ϖ�$��M��@�E���6/Y�ڜt����1p��܂�9�;���ɟ�F�9�ه[��/�{���U"�>�̓�J��ݹ�?]�������0@�.�	�{'�Sd��a���."ըଙF�u��=��H#���i��
�F(q�;~��U`�N;*4�B!���#��J�\b�k-k�`�'3*�tJ+	�|���4�D6<Ew�޾�ʩ�2�����zX�LA(���{�Zi�й@��S��ZZ����1�ڍ��ln�2�h�gE�4�;�7²����ě�@ΰ|�l�&F2�;��0Ũ������e�Y
z�a���N���׌Rx��e�7��C{K�����~�����[��lW�r���ަ�u�"J���6R����[�!ňzW�r�ۂ�Jf�\!��{�IqnSF���%���
�g��Ԏ'�S$Ct��Ӟ�Z�V����9컏����k03�>2Ǳ���JC�Y����U�S��(u2��w�z�u��D�u��{V�T�F������異� $�<�R_	�����2o�s��k�\�[,{@�}�h&l��G��v��Q���慣%vv�г+��Ъ.���B2���v���4"��ռ��*�*�-��Y=R�'�'<��Q$��� k:����^9cpnh�{t���P��gH��s~n��Zjk����">�R�f-)T�5ז����{��RL��"t}�PZh'ߑx��%����t�t��֣��9����f�0�E�"���|W wڌ* H��6�zF~)crz�A���Z:��ԢBc�@Se�U*n�K�nqrJV�;�bn��!EW�-X��s� B^l�[L Ϡ���v0�KI���je_0�@�j�0�����>z t��+�'�nA�75��Hq\��Bsrg�L9{��b\��s1���>�W@��j��Y7���4�L[��/�,���1������S��[@e{73[(���#׍�P���,ѝ����r`��k �^` �J纗�.�␽f)���<3٦^�u?�)I�V�0܎��	�jw@����n��hl�'ϡ����l����
�?ȧVD�D̑�)��jR��S Ԇ6����;�������]w��J�a� �/�����e�����C?X�3iڏ,��b��m��m��-Bbe��mF���D��"�z���f��Uzb7�̑HE"��C6��|���
�9��ʹ;)�aM�	�\	��c���q2u���ǩ��\A�����pWJ��ɧh�B���3&�kq�;��B�R�h��ybs MI6$cďeZ6�d{q����w��y4�u]� �!/�z$^���2��`��KA,=�mެZ���v��~u�&�aC{�Q�`X��o�'sE�^�N�I*�T��̔d�,�����EeQ˷mϏrd�fx�DZ@r���a{ ⼀��P����9-0��_���w�ћV1	��{��/�FeV7���vD�c��)>0%��t��1|�}���9QV�ah�ި��{��X�=��r����_	� �1)^�۾�lK����v��Nm�:��PL�ݫ��G��� U��҅�����&�N��� /������PQ-�S�����X���Z�F�Vtz\�+&���`Z��D�Z%:}�~o�q�[-n/���\�U���듯�1k����6���]�p�6M%"P۞��zP�u]���l_Y�G�(Zf3ȊA��Dn�$������F�a8�L��6�����@@��Gb���8�� K[O���k�����mma��?�Ej{�qH�^�@�qJ�L��k3I����K��?��TGa��Q~����Pd�'C���'�a����;�l���>�K+�aFL;�BT�&�}"Ix�d�b�vrP�܍�7}�e-��޳��l�\>��8t�ٙۑF;d� �#Ei�m2�8M�xi�G�g?��G�SJ�j�}@o8M&*p��	U�߳��O�,���#�D_L6��,r�LMC�.��'�"|��ƥ�3�nk^��N3�\5�trV�F��3&U�K�����2��d��-}`�=4A$�x��>e`�?S�|LX��4~ic���ʠ�r;�_fC$OvEG�f7h�bT*��7�p�<I�SDW7��Y�]u�'�����_5^�>��63n-ZKA���6o�\�Տ�ꕋ\q�����?�9졷G�@�-�V������p�@ܳ��a�����5��MXM]i�����{�pG�%��@"�E��¼�|a�^�4ǁG�ۜ���za�g�6������J�8�a�]͋����!��~U)f����ǁ�zF�u���IF֏b��+�Q�*vyp��BP�g!!���x��C8j�����m���M�ys��KRu��<����V�*��<åR��'c�_��x@���Y������>��@1 P����	l⿒��r�Y36����L�l)����t=����RA9��8x�F��xt�ÏO��s\��B�oe�].��"�=v8��(�m�=���"�P7ة������Tz�}���K��K�08�{ėnC��$���6y��H��J(lU)S�=}���lI~Κ�s� ��M�O��(�j��R�"�yX��E�t�w+��RW�)�:�B@y��:�����|;tY�"��+�s�()VχՌVM~G���i����Yh�hZ,	]��z�V�q�������A�&ßD�b�R�Gl��V����3���Y���������~�2��t���Wsr�3��%>L�����Ҷ�5�ڄfWM�:����+�����E�I?���]�7%ыg� �����n.����M�G2GEPo����װ ��Ϻ��vN4:��xXp�'?C�ۢ�!	�v�mZm��p��t���nH���2�3)�I�;�}�P��A�b�؏d{��z�0�3�	�(LE�������הϙW�eb��N׎�"�
-A:��C��S;aY5�Q玺E��ϫ�D�Q�ʕ�b�G�Ų����sp W@��E�A��>DV�PV��+  �~�*��Y[��v��lf����Tu��� �8��o{l���d��6��<��������a9����-�[�u#�k�y�J)��h�����GG5��g��m��9˅6�ʢ���5�e�6
D��25���0{J�u���cfQ��F�l���L�E��k��6�b,Y.�mI��;GO1���P�Z���o���!��7D����qne�m�" ,���7gƼ�TdO@sVL��r��A�c*/����#�ӛ��e���C�d�g0����M�9�z�=���Eo��1�7_A�0�zd�����Y�����\� ��ɗbߖK���v��{�X�{����i* ��Ig��0�ʳ�� jYr�#G�c*%���uLdg8)�c�.�j�nP�1Q�����^�+D�U&����9���ff:����K~��@t�-�cB'`�!��}�l����Z��?ӂ�n[
0�lE�R��^�����ulM���Ul�L�,�#&���zw��K���*[x�s�6�'�ڗ��)��1���0 ������Y����Oɨ"�#*��,�n!K����J"��pIʭ�T��M�NB�����X�Iל�MH���l�,���yV�%�f�_fA6G��(nC9��Q|��9�4�������Bny"�7��d�X�v7T�	!ǅ�|�7�\�
V �HLE�'c����mL���6��`��pMC��Cv��4k�����)h�V��#su���iF�����o?je��1tz��Eޣ�Un�����B#��s���C��m�3C������o^����R���Is�j��Dg@�ݥxco�zxS��1���2p5�&����fl��c��*3��e��`��%�V�y�Y��-~`����ݥaaވ��{0�-�m�2�s��i4��bafRn�R���~�̑�(���]%#?�x���7:W\�Lw�
Q��)@�1�������}�D��SfdndiL�T6S"������xl��C��� 9	I�Z��5;���������Wc�̞w�SA�|�}O較�q����Bkrh�8Z�Z���$(�ŀ_v%a�j*��f����X�r�����Q��@��vD	Y.JJ��=[��W�@̱��o����ح��߁�a��c��Cox~�G����_�Q��'O*�����^ϛ��1B(�3HU�s1�������0bɟsUYZ�5pK�Y�`���THe��%����J�]3nK^��lF�>+1+k~$Bǻ�"�f��]�9$�x��v%���k�.�gW����0khG2�_�e�>������4���{N��.m�t�mV�`���ˎ�v��5���Q�}.z@�c@տG����-��o��!�0��ΰ����X4���}��^�l�2�YZ�/^z�Q2:fP/3�y�|bK\�0:"<ekQ/<����;����z�@���!�'q2J� )�D� 0��b�bEG;Ϝ�Mr�l��S9���ݘ�1x��b���3kyu�4��ܔI�ޮ��Z�PY�8�w�FZ%Qds��gWזr���3m��5E�=�MB �5_�b$����
����{�O�o�8���":9}��^�����x�'�ֹ�U����;9�E�|�	�-��ӱ�m���0bJޟ��M��I��m5�Q�@[>�Lչ��t)�(W��MK�
�|�b�k�#�5$NF���Y��+�ê�����V���(&娵? �L�r�82m\97�T�_�5�G��_O�d�ڪI�x�wȑ�{��ww�y�D�j�ү#3R��0`���r�b��1��P�<�^U�-�5,�6�T���3^z�_�s����������������q��Z"��a�\c�v���Ï�9���Ce,��������廓=��Z^��:��2r1�w����9�,�4�Y��)��[��DNo���/���;����rU^���U�&���LԘ��uz�5�O��|����������D�9l�rS�na�$��U����ȼw�>Ĉ��/��88�71� 	BV'D�ml�{�"���q�_���@p!A����O�L�s��H�D�mm�]�����2N��D�Nص�f��-��6�sR��ԯS򦱇�};m��CO�*�0V�fw-�ո4.���e�ʆ��~7IK�.�oa�3xA��#��X��i��L�$����%�U����M�F�}֬��:�0���w�Oh!�q��=��H�*ouŹp�pTA*�'�h�*XJ�t��MĲs/�vw��`�U�*��u�P���ٙA}{ͯ	��(�_@���W�*�2f$}&K~�(7$�?�1���X���RW�ޡ��h�%��3U�c���]�6YN�N6a�o��-zE����B��_��f]o�t��E�����[%��5�����:��~/�	ce�t[�nĲ0ك9C�?�k�/��$I/e�5�10�B�7cx1��d���j�h��V��f�D7��.�'̽�/�U�}
Z����x��v��~��w�Q�U1�h�]���b���֮���Hz=�fvv�����]&���A�F}�we�7ģ���x@[
ju���F��/�h���P���V`8��cv~�SHM�[El|�/�#�ڮyR��Ɓ��H/?`�@p�1"�4)la�Lej�Q=,7_%P7&��Y0`9FW8t��W� ��6��qz`gl^qXB6���jI��y���(oI�P�HFU�4,�DjY��Xy�n)J���1��*m�J0$�N��k���Js�*�"�K�@��X(j��J�L���'˪�U���i�vY���=�k9�ޮ�Y�B���7o�&�j�?Wȣ�L�)c�� 	7��m�<�b�iʸƥ馊�n�l�o����I�:l����<s�����ST���~{C�<�=�z�Z1M�T]�Vh��y�*�ܼcwb���K�ZJ����臷D�ٌ�!Tqm/K���Q�H��]w�$%��JJ�o�@�W���j�E�k��%S
|�w)�mώ*ӯ7B�T�ݦ� �Z��0"��K�úT8N�����ݯنR�xH7�ᐃ����>���H���W: �d��E9~1��y��S�7�U ��V�R�ߙG#3�����ix����<3��D���K�.pEqLT�w��}�`�=����;���tP��Xf7��
aq�V�d�6�~� ��G�LDj^�*�a��^־
�^��vbr ��]�����) B����9<Q4����ja��Y.���kp��J�i&D{N�(Z����󴸜��ԅ�����ħ�A3�u���l1�r�{�~�V���d����`K�)����ˊ=,��u/*ۦ�7c��}Ŀ��%���J[k'd4^͹z$D)BQ�?���=�j��í���1 �
h�@�_����ϙ_ư�X#DP.=�S�9���O��n*:�z�DRQ��aL��]Oz>8�S�v2-ܹ�V�ۑZ��z�3���IB4`,ὢ�WA�~�,�$@ʣy�70,�h�E����'AV�|PG�diԅ���NE���G��V�g���[,��Ud���xN�~7���v�%���@�њ�����:��O��#����4k�0;V���ڔdپ��f�uC1����9��B��7>���-ʇ�JإC]7�4ء4VM��<�3�>��gejs��)W���D'kWb~���3#����oƻ�9Vt�m�l�S���F(�Lu�R��`�+�)������.�e-�Io��#apJ[�Ѫŝ[�ً���Ck��:��JJ6��K�����)�����/*���̯c����n�����:F��E��C0<k�1ssEdɀ/v�S�z���<8c�8�]-��s*�y^5�,��֓�o/9���(�r�fXP��'�	�k��睆	Ɂ�V!Qf�	����%�fGij�|��=C�8�>gG(�ނ�K�{�>��AYW ܉Ut�N��"�)�y���=[�3��Vc,���0*W�bI)�d9��:0@�x~�[�\�)���w���H�9R�~&���ϭ��47WO�L%ȴ�S�֋�E�Nx���j�\z� ��z�#L(���Cb�A3@~�\����jX��3���
Y��^2Z�ݷ�r⻖rR'`�
�
Oѩ,u3����i��n �u!��.mɎC��C��O�{��^����}ӟ��JݏmU_���-� ���4!B���u~�v��;��l�ågP8��e��m�Nq�� L����>d&cF"=�L��l�+�=��GD�=LH�=����o��M��P�%H�T�H�*�W��okfz���9�Ø#`�sD�4M�%q���l�蛡���.��^̏�1�u�u�`� Ή�<P`��dvv���߂L�
d��e����L��l���]�'WB(�x ^�deIP����X5�F�r���ƬP�hp��Ux�ҡH~�g��'�,���l�~�}�[��qB���a��Ҍ�S��X�nA���
�NR��O�R,�o_.́�I����ko��9�z�������xhUK{1�K!�j�	L!�̔��E:��:���̷(��c����0��)�_��s��炕77+��>R���"`)yj�li��.\4]��bN`%�-<��ןR3-&rl�Q��r�|s�v�F$&����{� ��P�o-=%�o��:�D��?��al�V�M�,�7�?��"T�-;4�a:S��>f\�g/m�!ڂ��5�XRav�%*"(��D�"�,�N.�DA���psd�ZmtBg��꿟3\kd��j�&[�p��m�+�^�N���<�:&D�饍�:�3�}�;U1����p�IC,	�Ū�Q{Η��K�϶B2cˏ�25�/���ʛ.�\	 �7&�M���$�r��!K���rbdнm�E&����n6�2F��4а2O����k@Pt�=#�N� �� ɶ��d3K�Ll��T��'p����u�8@Őb�㘩��'�y���a�����MGw�%�d��_�"�M��
;��Շ���P2S{[�D�����C��)� �2���(�R'�
�Bpv����!��"�.����?W!/"؉�=���1��:^~_�D�zх�<��;���п�jf�}�5�Fy�5��h��Z%�Y�G6���p,�'�	]P�> �}@�����>E�R�
���s���	�'�O��K��_�J���|_C<�BA�k�g���$�]���o2A��{�.ef�(�\Wo?+V�`������=8<��� �N���#�i&	 �v��7��?X�{��2p����Пr��k
r�(C��/myWjS�]Ɂ�������E�3\ؗ.O�^�I���Ѫ#|�N|3αq��ド������Z���Y�&6T��H�{�5z���R�/s��Y�q)�����}�����G�����nd�gN� �\�\5�]�L����#�r+�=�0�ݭ"�H]�m��2C`�C��d��S�(������0���Kz)~�+�_%]��WUc(/�.̤H��8�1C�gDn|��|�ΒQ=����FCu��G�w�9����� �<6^ h�S�r%��,��nI��eߞ�/�?%R�������X�~}�������~�9�8�H�7Ҹߍt����������k��J�ЎO^z���j�-��/f�J1�^R�{���(�-��W�
�/�ij��q`�9�7��!�h*�>��.��?���>	bE������ɝ�A��+I8_al'���]�q��׽f�N2g�[���}s������/����w����
��t(�j�n1�cd�{bg�CL�:�}S~B�2�?�&��ɿ��Uڏ1��� B"P����#�-W���,e���O�g��MȣyUo̦�)���6��)Y# �=�?2�p�߯"��s6�&�U�n�Y�n�z�L�[�Fq���;�xi�ǟ��l�&@s�?(��sST�9�q���n"*QX������*@��~ W���TKRn��2$�t^�����:n:@�0U�9])[�\�� �7w̞��y-��$���|�St2�Iw��^�KIG�&D���>}$�·�����-~��~�kRf��g�M�?<u�L�9�pع������z��F�]CpC]��ip<<U6�Ah<�W/s���?X��\!���D���&?땱�T�u�L|dd>W���l%'R�C�rפ���zBi�w��=
�\)Q�P��/�qnm|�����s
=�j�`�|���9���|���
�Uu!�B��χ)� ������Ɉ�q�#��}��I������ƪRc;Xί?��Ò����@顐c�n��)�=�~���n�nV�%b��.�TP�J���+m�/H�@.���fT
F��q�b"?#D}-�Y�+b��5�O�w���O� 87Z@b')��"����������Fr�,��f�(�q2����F?����sB��8���M����H��u�uƩv"��D�/�$jQ���	�m�2r��Ee;��!z��_o�̝�+$ꆽ^�-��Ը��\D؉�Q�S!�.�c*S	�z�]�4�o45���9���������[�k��F��dLv4���W�I�x�8d$�ĝ�"	nV��j65�tYavj��P��zA�_l&\�q鑶S�Q�d�lV�`L��l�;�UM|��N�>��ʐ�7���T�'���)b��C2`��Fu^�!��H]k_~a���FԁO��ڵ����c�'�-���7� 5��~v��q�M,���.����u�N�F�F�t���b�(,���Օ4�n�}V��_�^���W����`�D$M�^�Y��@1�r��y\�-7q��p��M3_�P���&��F�T�p+\��8,�C���?D���5�� M��	�*6Ұ(_���=H�"��X���I�ӿ�	�R�Oy���6U����T��kF�Ҽ�6ɘ,�}.��� �����X��N��3J�fU%�5/�@��,Db��c]�D#�e�0q~mCL&�;��'��Xp⢘��8cu��v$D���Y�J�x�C ��<��\9\�vUPU�r��5N1�~��[khs45]�9
�WlC�L�Zk�N.��j~���E�
b/�
�e�k�/CNӐU�������X�RwQ��
�/��3�$��uM쯕ogC�D��GOxK��E����p�N�&�-�$X�_0?���g�l�1~7�.��3�V1�H���ZBWv�������.L��
�З��J���~.�y@j���CQ�H�m	(�B\f���S�kA�-%c���}���Mi#�����T�Ts�{��L��yp%#��z��� ��ܨ��?�ė�m�h�m��@?�ݶd��+�ϫ՜m���M���_l/"B������~����X���S�] ��nK�t�L���������gn�Z�m�G�x�I��P|*�Ij!�
�	,�.%��x N�r}��?d�j&X�ej�dA����C�S7�#M�v��J�EfHN�!��0����3Ի��N~C\�jh�R��\�c�z�ͻQO�z L���7�SB����I�o�~M�g!e}����C"����G2QY{fwG�e=v��0�SfRT���āy�ʅR=ͮ�_w���
*����JB�U�\E��?��!������A��-���@w}`��Dn˛�'��`��h�4@��
~�<nQH��#7��)D|�B��{��{u�JD�\��;�q1��)Χ�'.7?��Ho�E8C�z;�T},��ۮ��$]�����>,Aшm��٩�8���$�C_��w�		 �;��pqM��.*�7�Q�LoH�^z[�+�	�~�as�JR:M�@�$O�C�_�YJ�f�:W�➚$��m�ك��Iz�D�S�B*����K4��J[<����e�u���.p�F;ЪGj�����#�#NeyE,�R��=��~h;H�P�PV�8���������N��<�R�U��:��T*�6,�V���CcS�0	�GTM�[�n�3!H����Ϫ�f�UYI_;������[�@�f�5�J���|����3�*�^���C�b{���5˭I�+T���"�r�>iiFϷ�+g�����q���FH�"]�Z�-��� 	&xs9x3wϦ��N8���oH�gA����ÆF�n���l���;/�Ix	�c������̏�w=�ƽ�� ��S�	Hcp�iq�of��7��\x�K��e���{W�ؙ䱔�oN
̣aIj��% �j�-\�����m�1*a����W�']��̴���2S��m/
gS-z峵�wb閉�(����I-A7�/J�=h9�Ndm��y�wh_�"��S�B��p�Vm{�����Iú ۻ�:�́��ԉ����v��m��o�IL~��=��<�s"���+Z�e�ZOi0���}tO�Dv/�� �ᇜ�$�j)�j�s�G��٩���NY�4w��3K	�p!U�.�@B)^E�Ξ� �"}�� �=� �嚳�Eu�&�rx��l0o�u����|s~b[>{=)��ݥ_�f,F���x�գ ~�Sweh�|t��,���K^�ا r}��wRpu��)M�t���٘>�(�+Q��!�����N�J�� 䧥p���ݭ��f.	DEf��fM��p��t�qe}NZo4���l1��O�����9H�aZ�𖡲����b{yA������3�Z�P"��\Q��	�֠;��nϊ�7H!y�I^)�{#B����ޖh��N�a��w�<���40|�B"��Lb�����fj� Xv������N���L�ǖ��fg7;"o�c퀒L�V#�V��U�ͪ���o�W5²@/cl:\p����2�bW��?�n]������:߈.���n-B���c7ٌlʜF���"~�YOs�֣������<C��>���&.�O��H����Þs �ye}.R6S��j	�����i²�g�&H��ǿ��*��3>��P��ڈ/>����G����%1a����N2M�c��<`X���:7�#v����J�:v��p�!U}� �GIw�����
t>}z�a��DUϝk�ؼ�.��Qz�i.�0���F/����1���:h3�ɤq��5��ѳ]V�q��������3t���JV�p�	W�K��6���S�f�_r��`�)Y�
��3&	%'��������*��$w�Ր���n�#|��_fĕ��y�#]����f�!&]4���:I�-w���Z�T��u7U������"[b���Y�����l���Y���.	vu��X;NK�LNv�Zg�$�A��ǭ{1�8`��X^�_代�E=�s-4K�e]�,V�-���5�v��m�!�}�x ���|}<�^�$���Q�&|����_�̸���w�+o��M@bqt�ߚ|�7\bDs�, �����Tnm�}�U��i�
EnoiTf̋C5՝��A�[˨���������gͼ \��f�Q���>�����c@As�1�<�H%o�bTV��SFNe�ņKCo�|�!��R������cy��t�F���KmRoT`�1����Y�j�bo���nx��wđkW����o�3�3&;5���� ''q�T�P@�M��8v�&��P�A�mʃ��I�90�M%��$/9:
��Q��zY1��$C@&�m;���RVE��:��p��5��\M��U#I�L9��Kc:�W!n����TC>'�4&t}�_�dr�Ag���wr�#��B�#�B Õ�K�r��d��X=Er����bܮ�Q`ߺ�J��5�^V�ͼ�lYg���VL8�%G�A�&
�<�Ea�C��g^O���-ow�+j��F�������W!	+Q�y��
;��S�	��V+��3,Knj���3��4�}�6x�+*Ϯ%#�#vl���.�i/}��N;��t�g������n6I�q�п���)�ON�iW�Ng����bis����S�_�]ڭ�|��ɋ"?6��S��7uE-��}u8��9oet���g�ǿ�M�b�X�L��i� of^s�W�5�ଜ@Q�7������B�M|m�:�Qe.3@�_c���[�'X�h����%�`�j�&j�J1O��js_z7��Y��U����!�?�7ȡK�"h��!$��jYy�mM[��VXػ�r�@�#]l)�WӇe��1x��0��������e��U�&�Q��ϸo�{�{��h�C���ZHz�䴚�'�� ��5��(��f�@�,�M͓@�!>�s^���i�r�D��x.��vs��@ے�+�?��nXN�*AM��Wі�,x��I�}�Yh8
r�����I�b;M�S�����h�; ��L�=�hd��
%ɎO���߽=���<��LK̴���K��?s&��>����u𼆝�K.o�q;2�/�<���]����>0�'������y�j�����Ug'����T��;�K{Acw2�Ռ�K��'B���C�����[o�m�b�S�� G ���=}~�4�^���n��p����/�*,,Z)i�������'��{�L�	��6�y���W��lo��{$>��k���b��W���X8�`��D,1e����s���#�Y5����H��e�HʫFv/-:�Z��,τau%�)�����D��S���C���j�Ux.���J?�g��c\��
kذ��=ړ�F�@�Ɩ(�d�p�AM-I��Q��7 H[d�%�E��,�uI�fP���B�U�9>�����`}R=��L�|5�%SO%m������[Hg��aw?N �$�)e^)3,a�t}�y�@�!��ĨTA��Be�ԟ�2X��?ς$B̆�k��52����غ?���ӯ@[��̧}g�������MR�7�f��I;ܔYo�}j�]�@�P���^��u�����[_�:߶��x꩚~�[|l*�j&x��LѓFxA�L��^�`C<���|�����g�¾r.;O�%��Q ��+B*���C���Q�E���v!۞��:7��Si4���5?�i^�+��쏕���X����*�UV���P U
ػ��7�k 7��4 mS&H=�8x��ُ���8�a�_+�HO�+��L���u_RZY��f����R��x�W}���i�ʇ���A�6ԡ`�)]��WږV�*�ǮKU^iMI��\��E$��AQ��u�E[���D9��w��Z�3]L�]9�k�*;�dG�9��爐�;�}�yU��.j���v����Y�aj���Ϳ�1���쟡b��CDj�g��S�������W�r�qN��1Ĥ-�H�S^�?��|�~����f4R���D�uݐ{��A�Yi����)G��[r�(��b`v#��_�M�E���*��#|}�a���4`&��z�`���>al�!�[e_�
�8�
\�Ǖ;������`.!D�p�j�i8ڇ�XwÄJ�t�Ɗ�p�/r�Ԯl�@f�3����BD��]��Գ�Q/�GAB�ћ�I`u�{{���w2TS�`Z�xv*`8!7���9��U���� ���7iSӀcb�=�A���!����J��+hy<��*W>���. ��S��p��;�>�� s 8�㾬ַ��m8z|Y��)��I��p<D%�����|u�y���"�.+��6���S��6�_�Z�4ёB�ҎKi�X��!mkwM
�Է���V�C�Yܒ3��K6�^bX�ɴ*���Q��!xW׸o k�,���~ �_Bvl,t��NB����GAS������.wNąR݇샨�[�6I���\�L� ��[����l�-Y� �1L����	�����2Sሂ`oO j��W�m�4ͽ��3�	&�0�ߢ#�7�fMG��(�딕z*k��s�6A����>)#Z�6U��f����h�(�M�3:��&�9��^
�vWnL1m3�܂'&���u۸�vkltN�s>�mN��gFu��;�Hce:��K[6��=�,4���3�V����,|����M�]KW�B��\oZ�>=�{��r����ܢ�.��f=Ԭ�}IK��������F^:0S�

~�6}�p[7_�yja�0i�΢L�A�_PIK���,�_QFh75+\�X[@�{�k���>�0N*�1�+�M����ކ�i �w���`�ǿ
 hB?CGQf�T�r�x�"��@}D�Ţ^Xwv9%�)�j�*���ؚđd��F�wDL�Z���z���Ĺ��2�D�����:��ګ�R��BbN�8�����Bg��v�j9γ���yj]P�@�oo�J߇
F����L7�#�)zC5[�qY8a�*>48��_�S�"��ɉj�(��t�z���8U������n��.,+��-#��<�&�sf\D=���j�����A��,,#���C6/9ɤ��	�ր�0�l5��Ŀ������d�)�lֹ�Q��@��tY��w���e`	��vf��K��g�@�	��"�]����֚�� ��-^�j��$}{j0��D��睅
@���Y������#��C��L��å/� �(��.(j�lt��:ol�I	�[Jpn?��gҥ�wz��q�G�����(5!̰�4|*b(Uw6�,b�V����&�h����%0;?�~D1�D�b@�Z4��JUʟ�/�F֫I�l.�l������A�~���{��F�l �SJ�O�M	h�nd'Wd���V��D�1th�����v�Dd]���`��b�e(��paJ����t�80��Z��	���}�Jq����"��������#�]{+��U��Q��>HZo��P���>�� �����Wp,����(����p�Mz1T�^g���N��}i��_yXS���[إ�oT�1������I�l���J���E�/`����CzP�
Փ
K`4H�
��Ρp���Bl#e8��5���&e��@�V��g,�2��G؃ݙ��Ym������0�(��r��
)gduC�k毱$�@��@ELnm�����?V���E��y�09b��
I\�zP��Q�bO#��)��%%�PE���i���ڕ����m1W�7#����p_8&0��VÕL�`�bL����e�Sly�~93�5J�>����i�:�ij||V^��UO�V
�,E����X���X*p>y�w�A>�Ua���a�FU�l�2��{�*pG�b�,3bxQIwz�D�ȉ�K�fU�Og�RM"N��+�� !�M}��@�ǿfH��29�?q҉�׌�W����xӟ��*���I�nϺ��S8�Q¬�0$6�V�#l��� �����O(�vo����_U�z�΀��������c���b����	��_<f�}��@�h��sz[~�Q��!��[�(��СI,4�d@l/H5��ǖ�1�t���T}-ޒ$AY��I���M�)<r��&=�j׊�P���v�IF��q��G5�2��M{�~��D=!{}J��)7�;Kൾܟ�W�p�9O|�&����%��m��/b�W���`���ɹji���ջ����*���1� ���s�-/���B䋖�L�l���� �����nDЄ���#�i��N	�o�+\�gH�TB�rw�&n.���r�u���c��m�����M/��E�v�!��zqr�㒰�ق��;6d���Uo�R8������H޶0b�+xj����-�v��R�i��E�v�gzx���U(�ܕ��n���d���J�n��sm�y8T���,q2��[��ǀ�T;�
X.7m����+qC����'�U������/��Hjs��|8s?�`ze�h�l��K�]/T���Kv3�rsR�
G��e�,-�"��Z�$�ֆ�!І� ��H��X�U-�y�ά3�E�F<m:.}5���l[ڕ��kH��\�N	sG��,�߹ȯv��=4�)?��=�kJ�]zq=� �j�ւT��D��?{�j3��Z^
�ca;-��enp!J������`7���c��/v�[�U}ȁM>摲w"֋Ñ��q�D^r޿���3.�b��$B��a��� ��\��Z�-mY�2[ձ)/������ �e?�h����	vv��	�i�wnb�O<��(#��pޱ���xu?8�iПz�tB��Cd\#A,-_�}�BP����]tU	p�"[�G��)�S�9�NB9��"�̷��,�jZ�z�".{�+���
��ˋ��Z��~��^����dm��R1�h˅�ֵO�9�rOM`Yނ�8�O�6�0 ����b3�EC����׵I����sSҲ���xv	�r���pY|�-����,��1~�ҥ�6p-N���Ѭ
"19�^��X�jH޿sr�k��?c����*�����F�.h�_������T�6���H3�M��`�p8y������zX2����>�"��m]l�Dtu��h$�����MG���VE)҄l%^mN	MdOWW�K��N���y$������9�ք�#��:���Z��Vf��+�yƑ�-o�io|���v�3ǎW����T�?u㧕s�a�珧m$���3g�.V��P㠡Ԥ�q��t�0���o'=�l�-;��)o��^�7�<�!<?�Η��q�?����lG�4���w@Gzi���wh�����=�}m��TD7�l�� PU����u�=^��ۼ��5��=f���d˼�('�t�{��'+u�8D!�We�D trl'+�S&y0���WuM��W��c�h;@<�apք�gd�褆8]��~d��H<`��Ґ�)l*��-�P�	 t��m�'�w�C����KK
��/�wT��UwF�S}�&��Ngem��=}��A!f�R��v%�&�6����ڍ�zؗ<uf&������Y��#jP���lz���[���g`؝I��f��/����FU`3SHܫ��T�����>��r$�A�dw�Xy_���x@�g��rd['�eȧ��즰�<�0=�/@\�)�C��[h?���%�4���y��-���������A�9��K�wҖ!T��+:HaE�2]D��9�I��E�[��#�x��J�����͍b��� �F��A�FD@�+��D�u�C1oQdU{D��1���ht:�+yѩ�c9��C�Q(��>'ز��.[QW���(fch���R]*I�ۄ�ۮ��2]��-+�8�#�\���k6+zJ�:���Br>By��o�F;���L79
5-�6H����C��3�����qaI�,���������آ=�?Jtub�]/z���(/��h�酮	�|��tK���+9�w���F�%$`� ���]�o	}���upr����JFh��������S>d���Dz�����Qc���s!�+ �;A ��(Ias�MV�g߼��V>[a_g�����Dx^�p��:��&?�����yV�@��V-���b�!y���M0.�:í��26`Ah����Z���DR��P�k��=o��v��u��0��]{Ӳ܋9)��T���%(/=>Ӽ�L�c�� ��a��W���^&�fq�1B�3��z矹\��p��A.����.7W�sB�o\��]e�o�ū�1`���O�p�.@�sP��쑿ąl3�"����_�r�Bؘ·��x?B�ק�\͔j/[;�����q�<ľ���-y��q�[�����RM�ɏ�F�JXS��S�.L9���#���8j�d�$�y��zq>l�t��˿=��ǣT�$�I�F�[{�i�
�����^�W��n[�����_���ÿT���⦾K��d{}
B�'!|DF���L�z��wp|ǜ<.��7F��;m����������v�a��+��6�G�`:��h�xەn�]�/bBƠ����΃)�;���0�'�e%~�'4>�~5fR^�aR����6I;a�M�UB��.�}��/��f�?h���tXͶ�w�/Gǧ˂��_�a"
�D��f�w�� ������*���@��g>�2��� ���Ņ��#����(o)�J�,;�	%)F7d�?&���FL�WZ�H�� ��~>����s���g�FM�p^�-M+o�7�&��si������{�y����{��3J��S�ԧ���(ńg]Zv����6�8]�)E.�؆���*@��MknV�,��W���Լ�,�F_"t{-`å2�tI8$���E���*<�2|h�v���Y� ��B�;��:~o��ZY�D`eQA�@��*�0���R@Hc��O\@�;M��k��������4������o2E}M2 ~eW��tN�vTA'22ΜbT�겘:95a�3P�~���H��
~�����M:{��@u�2�q�9]�sRZM]��!��c����[g�Yݔ'��DLQ+�r��x��B��z8�������H����ˏ-a\��Ly��ݼ���H����;u�p��TD���S�&�����-�my�Ra�����u� �xk٬���3f�E�N�ԫs؏[9�$�~�Ym(�o�%3�No|.	��b�yn�+� ��%.��AW���<�	�#'�}��vk���4p�����l1��o�����6�#���	:��ګ��`�j�� lަ��������V�E����oh��.�y��,�?{���y����^d���Z3���h�}M#VX��k_�
�Lz%� ���h�{?��_^X'P�hw�A��>�Z�Ε��HM0Kg�!ikE��m�я�NĹ��+���ܢe�7�z)�7�t�͖�[9�y:m��s3���Ͷ:�F	���/1�����i6��ڵ�"L�C��Ϳ�#����$�8G�#	��DT�^7m�#=�Z@��@x(�]ye��S&.��K�G���*ռ7Dn��{SL_���ɷ�̑gL���0�٩��D��W������%�
,����_���4皶��(d��@ВR�]e�y�����*�Ȗ��|�O?��bz6ﴯAC�_�;��E��?K�0�1e�����U�Jc�?Wl�(��z�F!��x��W�!��:���׊A�"n*�*�R��q{�jT#����$��0���޹�cO5��8��5�W =4��)�]N��z/�t9 �t�O2`$Ú� ���ƤZdY�ֽk�s1[��]�_���7C4J�B��LLo������$eו��z���6��O�E��&yHo���G}&=4WX��1�գlzs�J/;=�V��|s���Q�$�q�J���L�	1{�.Lu��V9}�S��)|S������#�t��IO��b���hLr�����R+2��5�~2m~�)�3�����u�0�WnL4�B�M?Ջ
��\��3r��Z��Ǫf�E��������zR&��m��������v�{�3�G�AF��+������L$j��u�B�c7��]g߂�����t��߳Hڲa�O�B��b�4N���Fq�n���҃�5�%�	�L9���m�a����������%�pi�����?&zy5(>RÞ��%iSZ��ގ;��&�K����c����V�e����m�)�g�ى���-U5
M���)0�]�V�,6%Y,��
W�J��K�ABy�~Y�Y����w�	tM&C�����I:�b����0�'�Mm��nt�a9e�s��l8�k��N��k ���� ��� ��w�Y�<�6T�C���of��K�GWJ�gsA�����H���t��U��!���LZ�Q3x�-f&�j�X��z��6�$ӫU)��_�[�)8_���j��ʏ�>O��R����7�NZB[����&^	�&d�tY�X�� ��6օT.O6W��Mj�h�|$��h���p��M��)uCZ��F�/�p��]*�3c��'�ذV�Ya3G�
|�%�@�S_	W�WO�6�H��H�$
�o�����c,P���?Iۡ�h`1 ��N��Y�L��z�n�=϶ńW���C�.������N���M3�
[w�4�3�Ɍ)H�7zb�ĕ�q����N&�����φ�� �o�wM!��b��R�2�q	g$���#w�-B��}\��J�U�X��$;��K.���q��
��8VC�Vf�����*P�8/�y�oـ���0�u��*��u�Kt��}H%�PZ���~����r���u�2�h&�ʳ�����]'�qz����H]���:�����PC�h�����;I�r�jd��IOѠ-w�x���c���
��>Q�����(���;䄽=�#���q7�禵��
�Z���U���P�]U���[y��|Nr����x3��-�����g��7k�.o�Ҙ1��;Ih���\_0�hH�I�W�yS\N88E���z�[�R��SN�ʰ���1]�o�fMٕ��qޔ�J5��ւ��렏#N��#t�9�h&��ڪ�g�������	���D[���S��F�#�c�*�N�wl���r����Z�\"9��9� b)B�:!�x6�G�ր��M��VL��6��ۣ���E�MqkA+/�^O:W��6���c�:;I\s2mp�p���ŇM�)KY��:9�/��3w �#����(;�O����D�Iw���ÙH�U�
s������v��Ik*CJ7}�xhx�y_��GKob�{�4i�!�PW��~�>@����� �ވ�X������y�xs�	U��<�w��ʺ^ @�8*L�g��Z�-1��=���1�j�UY �֪��jc�3�����Ds�w�l|AM��G<�.�@��g��A�Y)��o�g�](X��s���kg��ٽ�'Y%{Io���&Ƞ0��} �|\A�b�2� �aF�	<�]�aJ��֛))]bs_��ʅ=#��|�*�ٗ�� aN3s7�E�|�V$#�(�?���T�H�&�2���P&;��s��[�Ǔ��80	t�z��#�pQ�՘���g�s!D\f��id�I*q���D9ȡ� v^�(�Q��A�P��Y����p��S5�b
4��Dpnz©�!{��*t�_,�pTc��Dc������8�Ǝ��.��`��[U��J��zv��9�T��B',�j�x-_�ȑy�i���"̒ ����n�1�O������v�E1�à�%C�$�2��B��� {N��!���utؑ>c����l�߰@:z�h],�:x�Ԃt���|@N���QLr���;����2��w
�+�W�=;�>����:2&�U'��'�U�v��v-�]>J���q�q(����WXCa�}�8�|�5t��_��9TϧFš↼����D~���&�7dH�S(�t+��E&=��	�=
R���b1��t~U\�$8����_��rgUR3�H�Wr����~���ũt5@�+w����'v4C�r,,yu���(��Q��>�)wy������pЇ���cI�O�x�%BT�Q۬�L��$X@ᔊ_����2.JAp��=�`,u��ͻ��J(�����?1}z���S6��5�(v"V�R�=���r�qku���xΖ�?����U����7ګo��dx��cL��/:Y�Pב���f��Yz��k]9�J�E�\}Ŏ��F�����[��03+�_ۻ�=�@OPi�[�����ԅF�"���������Y�෺���A �ʟ@0껇��-�u(����	D�ךW��X�? �~זz�v�����+lb%M�[{�u9��u�G�}qr���G�\e\#��R�E�4�:g��Z;e�J~��15�lO`=�F�d��Qx���4
?��d=�������u`���6������\J�z������z��K�������ri�����,l
�`_�=h��m1+)S��w��ݑ�.?2��)��k֎��g�Q�D)3���\�j[S1n�H���1�w#��?S[��7g��0���U�׿/d�5��e3����7���w_u�aXI���ǡ��ዻM�%-�T,�5tm�b�i��A	����Hh�n
��������m�"���aR��'��3�x��O��ʭ��U#�q�����mL���n`�Xxg_�-V�z+z���R�.D�04����@|P;�e�3B_�^2@�d5q���l-����^M�
?��Tf��?���dU��@��0��^�K�#5c�d,�7��Q��sdC#j��~�E�������r�JFb�%&�Mp������`��;�cT�ˢȁSWd��\\7��rV	+�}rT� ��c���'�c[��#�$��9����A{E��Ǆ� �O��s@47�r̂�:Mb���V-����c���/���:䘛�3M w="k��*(�w�`^�����\����#�#wG�_���²c$���Qٞ􉚠���R�K�SC�}���{Zq#��8�ºB9W�w�A��
������gL\�b��9f�{鰐��Qb,���ª�]VY����7�h���O�����gr����RG#Hi_4�M5�E�c.�ݥ��{��\��_�8l�jC%���D�k�hh7���y�ϲ����t���beRH��&�L�������.w6�ali{VlD���[ӄz3��>��ڟ��0�A`���C��;���2'����d�.���ȢD�M��l�4-����X��0_���AB���
.�H� 7�FoՂ�q������9� I�ŠO�mvELS�n�Ѐ�*o�}�!��=�o�AK���h�=,����M4��x�N]�Ć�2�#S|�$�%kC��1�`2{�Ӱ�*�S�~���U�sU�ZC/2Z潥�,0E3����ڇX8K�j?�|�gKM�BE3	�Ei� ��Zk�;w���r'hFmx�ȗ4~q�)M*��z��[�oհX�H�'G�`wvSGK�S
�b�5G=�-�~��_��4���K�ǎ�j�D����osOw{B`ͦ�x�c��l���ƜK��n��"5�MIg˄b���?�=�'3e���:!��������e��L["������Dm+v� k@7����hɁ4�'�r�k�4���R���>�W��ҝ�q��4��P�' \�7<���h2��weÞ|{��\l���9��,��X���~"��cp]{�G��ж�8 �����xHn��f_Fy���|"�Å�s��\N/�[=�K�G��v���o�k�J�PlwyQ!�5�d�}�����gd�ʄ2��;�����Ќ#��mGk�����÷��yf�)�7��l.�5�+���@6�,]�����2DV�����˳��QDS׫M�~�N;�R�l,��*�q,��d���B]���9:{���נ��:��6 �<�u��I��h}o�cA{e�ً��%k9fD"��+7$h ��\Vtl�<�&ԟ�
��kS��Hϳ�7-]��)��ɦ�Y2	��~.�4�w�C����)ks#����P�j�D��*cM=*�C��r���[W��5�xWC���F�������{_k�v�\�A�Ro��E���h7�pv�i�X�;[�WK�_�qKCt�z�y���`e�Y&]�)��s���Vh�*T�`�L	�����Y�뵢���z�Qu$���j�SLEΆ+�Qk	C�N��6%��]]�/����H3�>!b-<���R@l\������45bH�"�p�掻�~����/�o%~�y-N�V`|T|�g���k�x���y��#���z���_O�Q�!���^>�{v/^�f�%q5?�E�͈QQ+�Y�V�E7d���Pu�}Ns�j43sK4?�ñ�.:z�"�P��z80�
%���/�RlrYe�|bo�8�>��R��N�9��45%?P�Bw�����-$=&���!��;͵�oJ�	 B���a�3�WN�c$�����D&�ϰ�v;�����{��k��Q�LP�ᓟ&�㍵��(~0e@P��Y;�����4���� ߞ��[�� Q<� �T)��%gq�*�a�G2���^<ftW?�,�����E1kW�sf��^ơ���j2�:��r�����-9-1p H�͒��m�ǠqA5�c�6�7�h�j�[1�F5r��H+�~x�(��]����^��z�d��-�i��]hBF`��Z��<v���}6<���ş`Ԋ��Pv�]d�QQ�X��S���ɷe��� "Pu������4�^̦�lΞ��rN�u<頵̄D]�'�ANA�.���^?Vm�2���9YN�=�`g�8��_�4v��	س�`�Gm*A�_�ᔊj:P����W�/6�����̍��o���������6g�&w
�X�jsBCe��x�r�S"�O8D��}ȴ�um�)D-���� �	P�:��(R�teE�z3�:�-\Pѫ�n��@+C<A��8*=EùIl�Gx��;����f�i���d˕�g�8�n�$�#�K<A6��f�@�FQ�Ѡh$gZ�Y���ϣB�ۤ *����@i9��'�1�:��⧝����?�s�B�,�n���+�8��{��0�ĩkTg�)����A��I�X�����V۬�U��.&��\o{��(_�wޢ���{�b�����Rk֥C�-�ߴ�MV@7���!#��
�'/8�2A�3�j���B��40�/���v��Sy�W�\���Sy�r�у6�<X[,o��p*�T�7��M�\GtBv��b���S�r����9��]��8�O2��Iܪ�Xd��*Z����b֤)ӸmX��J�R����{с��s�`���T+��
��C�m��Lf���(k�r�^KG7;� �G����	�n�$i�Ƴ	�vB^����Ŝ���B+��4ѓ�)m[��6�3��/ӄ�,�J #SBn*&����N.����`������s}�稚.M"���g
�+��T���2�wg#F$�Ҧ�|��K�D^���y;�`]u��	���ӳ ��9�'�����R����C�l��&���1i5ǫ�xG"Q�L��H �g�J�`ĴB�6-8x�f�G EwA�I�?L��Ё-�H�Z�O�=�p
�.3R�&��g�|C�dK�5��ί�ѷ��o�Τ��&�(iX���u�i�a�F�
?\AA���fՙ��sQ�	Kg�M7J���)sr]~x4JY��1i.ӫ<�� ��uM"2LH�����
C'wfVt��mO7Y�,߃�l��F��LQafᯰ�>@=Ȣ"b$1IK�c�N�K�%�c�O����3�9�/d���
�T>�e�Y;L���OJJzK5,��F4�5�q�AƝ��a��Z�H�C����R�����>\��|.�
�!jU�w_�?ߦ���d�~f�����������"9%�zõ8���..�<�u���0�F�'�&�0�L�/��^��Y�P$h7���&���vwv�Q����QaR�����T�c���]*T8��-��j�e���8�1��[ٛ��Fð=�=�{02ǐ*�0�J �t2��(�0�,<8��?��� m��!�?`�i��V9���b��_NO�2k[�N!Qlp���K&�tz:8�nDN�`]��h9�m�Bv���'a;�����������c��ˏ�^<$���d�/wg�̼"PoE��q}���}���R�C3~8]R�i�?T�|����nQHS6��?aXB�Ed@G�Ä�Aj��Ten~�x,��U�����5���0��i\��g����*4m������R���)�äBJ���te�I ޿��!� *FO�� ��ޫ�ku9�g<[�����I[�RD��9��;�Hjl&��4Zd��G�Z���2>YG�c�X�6�e���@ �畨��g����%��"����m��� �b�:��j��Յ(*�kEO�.��M�1$��e�MC{�o�s�����y��#���Ɏ�O���hیF)�V���١X���b��^t�_ILゔ�N�}:e���od.k��W��4<_
dJpb�іá�Z��i�ƶ#���"ʇ�8�i���\�2�HN>�1��E��d3���Do�.ь4����6���G�`�=��-nyÇ�Fy��*r�D^�Ҟp��+���$L���n�Kh���� ���:�T�ɌX����;���G�O�f�%��s`�i����G8���h9Kh��P�o���3�1���^��"ʐ$�h�b(�b"�۾wd�!|�^"ԕ&����$��ۀ!p��`��f��1-��e<Zf!����u#[��h�w�9ag���r����
N��Bf�����FY&73���н`%���ee�! w�����MS�d"�S|S�d;4��9.2������Q�<j�#�`	�M�p�����͸vr؄���!��E�������O,��9Qֿ��q�^��+$`ȱ��� �9p���%<,�"������zo=�c<���d1��1G�}3�Ӭ�F�Ŏj7$�u��E������މ��H���������O�����ǻ��n�����{H��N�ë�/��Y��#e���Z%�ܵH�K�Ҋ����iaF�G����}Z��*�^(�P�����J�ںMJ�����H)04b䡱B"��OW��3Ǵ����,��U�e��@�bY���P&!o/S��W"�
�/`�(9�O~4�%qi�E}3	��՘;+wl��e�6�ʬ~\��DX�+_�I	%��~�犻�o{�q����pQ��K<�.bV咎�3U�
(vUO��*L�%���g��V��8_fϡs<���_P+��c�et2����'�Ta&�߷�sKr9l��u:��;J�$P 1�Å}��W�eŎzsϗ���z: ?�nyI�@���w� S�W&���W�X8��9��ad���oɈ������q|e6�X��G#�!��}6��ܬ��b�D[!�&�_	Η�R�e]�oR^5<V�.մ
���Co��r�w�5�܃�y��#�t%c�@���Q�冯Sn������&'���ER���lEXa�_`0���F���]v���ׅ�� �9/��}9�p�4����\r�c����։�5��\�h�-O4��3}Ρ�̾nG�jR�O�=����6�g��=��
[�(͔����qb�5M���@�E��w���
������[��\9��*�aI�5|�9ഝ����7 J��,�#�4�?գ���K&�@���7��fe�\��L6����)���&��q��"�[��"0&�SΠ`p�O�T[�p)�H���g$�CG��F��s�O���G �{��ZRz0��Ԩw,��4���C�H��_���gTs�<�q��f�g�e�X�ą_������ثV���B,_p}����I)f��>�d�WV8���_YwG*3����wO.�H���
���m8������>5<K=6<���sܥqͯmdD�^rB��x�)��O;�k�Qv�4/
#����C/���
��s��}�ٜ�V���u�O����bs���L̐{�L��i@+�Sb���A�b�ıF횄:
b��K.��ε�� �,d7��S4N����D=������o
m�y������#�\_���\i�_���F=���^�Um
�Q�V���mN>�/H�ܒ�5M`Y��B2ۙ�*^�*ǚy�q��w}$ɘ�aT�g��89��w
���nO��d�e�3�'<���n�Y+f�
﷼��Z�w�2��*) ����+��U
��2c^YD�Ş����h�'��ѱ�^�gYJ3*�0�k\ 1�}Vo�x�1�>oTa�ΰn�~3�9�=���J�������)*�A�r6HG�ʹh(o��ɪU�Ds(�җ�.�;5�i��V����y8���c�ST��&d��y�#���$jO����
W�"�q���^��gF'EQS�������Ǘ����0�i��x ۷�!��.�SO�ѡh��%�m`��r)�I�'�(�ݹ�uL`�`V.���v��V�`i�%hj��,Q�)	j�H�yL�������7��Z�n���n�σ�]�5F�t��3��[uW[YElv~u���F
1՗�2�bXWY�3�Dmk������{���Qq<�V������4>�^�e��~��lG����u}�J�ُf�������C�9��H�#!�ȇ�/�N�39cC��T� �:as�8)��4쏚.u�D�: u���a�nC�M��Eu;�J�z�Rf���=�:���1��
�vC�����ߎs�,D֒u�V �N��7ֺ���O~��3bO_��[������R ��dtaROƖ��!��9���<�2.;�>�/<��iX�؜\ʃ�CAO���aք8#� L\�;���)���vQ%
p3��A6�NDuy�L���~���8`�Z*+�����UU��0_��y(���^���;�����"T�/��H�R���_bXtP�V�U�T�bbʸ�I@�&y{��Q�4�H�=�Ww��JuWe^*��G1�C�"�+l��/�,Ե9���V�:�'�ײ��p��r�G
p��5�/Rk��I\0�#�S��6׶?Fs��\-�,�QzR�ԇg���x�SylrG�� �|�K�?�B6vC#\��>B���H�5�EJ��s�@"vN[d.�SȻF��7R˙�J-[���A�ñiE���/�"�1 ��jO��qƶP�Dd��l��M��L�vr�Q��7	�L<Q:��R��Nީ��1�[��H-}��srS�;\��IL_ʺ)l��)�L��$���!K�6 ���YE�]zިM8t%I�I9#�6�f��*F��|鮴ro *B�(�I��=�,����C����s	i=��5;��#7����K� N��!�>���:�|΋*���P��i�Dgo�}M������x�BAf��c�%ػ]�YGx��oi���ϔ���C��0"վlFfx����3���D� �z� *���{���i�%���z��h��n��)^�M��$�փE<��늕<g0��I���c�Olf+���%�њ�V�i~�����\>�2<�!� _ll����KU�����$��~'�x�N�C�-��z$G!c|ZC���\��}9�g�>
i �~���\�l�4+k�2��f�\:zֹߍ�h�yrW�u����2B��Y���Kq�NM����/�`�Z��(\5�3�4en��3E�'O�6D��n�"05'��L���ʾ'*x�D=)M����NϠ�����Z�?��������Go���ı��J���>�4$ �H m�ٚIr�[���e��Њ���1����<�\9���xZDhW��#��#�Z�=�D��?��J���	�q����Bȯ���� ��uQ�}2B99nKG2��c7^N�s�Q`�~����=�_�.i��:-/M\���;4��ё�ݣ%9�e>v&�:���������âۥOCإ������٠�2�+.�dZ����7�Y��i��9������/�g��
�h����[f;ǣ��|}�2�BQJ7�mg|��
 4�&9�O����+I�U3*~WF�v��q)�U��@qRL qu(w�g��׃G�
\�H9r��}��7��	�teP���,�h\�����O�T�{woz�$M7��D�K:�����~��J�
U�ǲa�.E���K,O��jl@��,H�fQ��m_S[���.̂���5�!źV-��G����	��q��΍��?;
B��?"����8A7<���C�`\m��ܽ�(W-��؋v��W�m��w�
g�G<M�Ľ ��#wu3���E�8k��;���J�" }�.x��	�J���4�8ZWWl���܉[�I�8���F�X�\4MdNޓ/�����M�v#Q(b�+T��?�'�����7��~e�������H&�m�ǤҊ3e\�,3��2]F���4h�um~�Te��02�75V������=+�%��(Q�d\s�ڬ�L�W+Z螾�mg�c��ـ�����z���w���9/�
ߴ����I���p�@�+/֐�U���H(�ʻ��Y��I/>�P��4��7&!���E����5����u��E�Q���f��rJ��8���0�3�3܃A�2����G��#������{>L�7�Fj|� ��y����ň`�Vb{:�?��s�-�	���"8�U�.��c�&Vn U�v�:&vg>�b'%�T�C�2�}�q���G�a����3Z�C6DmI���Kf���M��z����N��%�cE������	�L����,��]p�
&�mZ�v3p	l�hY�t8tw�·n�uGE���G0gO`�����M�9 ߚZ*��˹��/X�'��S%X�C7:g�y����/��zF�>'��N���#]콅�{L�	�*bC7cvxFi����cHیS����׬��^���<�i��K���=VE���n��i��	=l��u��� (�\�qm�j8w�cS���z~tqO�#z1��\	`�Pk��ЖV�?O�<��'�f��Ai����9>���gD#F����wn����W�Q��倣}I?� ��;���y�rF�J��t9�����ժ���`�9�53U[��#�HS=/��ծ�}V��w�-�'ԇ�u^߿c�
/����;\��sBNf*�E�����A ���.#~�+��O"y�;��iJ�d�:�s�a��}5w�|��<]$�s@vf�$o^'&�S�T�K �ݓ>_�d'S�H���Pg�sQ܇@�����%jC���-`&8���^'�y�X�y����jֱ�D�Q#9uu��F�;���JM~�j����/5U=�k����M��3m�:�`<��#��������rI�@���8��)IpIuH�7�di�`���iG�������g��Y�X�K1��3ߒ����^�@����Z����曟ۨB��-�T�H��T�L'�e @40�݋�VT�Q���jb��U!̫4�Dkӫh���1�Tن�I�@C����ݭz'���tҞ����y�BžJ�&(�*���h{:���!���̬�i��XM�r�,�rl�|.i���_�(�6}x��S���,��4U5���gUUF�t���x�ֱ}�~�p`�5C3+��ay�3t���$7���9h�H!ڊ�7xJ+�p�qr�v������xJ�`8%'`��,X�ELP��4����{H-�U8�1@t134C�#�IT��ؿ1d$����'���KUN9m�d�ۛRB���@)�`%A��=��q?EO��HRq�8S��(U<u��["�ׇwݐ4 ?ļ��Z�����M*�CQ����F��u�E���n33)ks�G�SO�m�뭚$�<�Ť���N�kp[�v�[���o���+p��2T"V�=[���v���:��B!�j!Em��I���Xn(,um���|N%�Eh8��;+�W���Ѩ��L����'ӱ���&�������ǵ>�#fg����m�V�~Z�r
ђ$��#�1~��Qfo���τG�K���~Q^��{��ϳ��W_7�H��+YYFU�(&�p�:p�}�+��i4l$�@�HWrL�֏Z�Նg��Al�֢"�leD�i�Rf��ݛit[�0ɫ�*2gT�����=B��ݩ��8�7 U���E]�3 �D���R�[0/�B`Ẍ,kt�Ď���ܻZ�\Z#-n�[u->r�CS��z��V���j�3<ABԪ�g4L��=�δ����\���,}����%��X!֪�a2 ���S�8M%�:'\r���+�bNz�}K�-TBSH��g,��EW�1��	�I:A�;��'�Gʇ^�xhHP�1f�H�����7�<J�C����f���޸�����P��hT�(P)oַ5D���-�q���
� N�U�x��v;c�N�Ōϴ!�M�&-R��cP�|�f� Πw�����Y�g���xX�An9D�aXV�QY-�®+�¹��S:��K��D���o��~���o�d��-�/I\��M�ř�&a��Js3gq�H�+?�`l"��5}*���?i.��:�"NY�wĐ:�	#�Un�JQlm$pe�ү
�'Dk��1On8k�����5y�1s�Ȟ0Tĕ`q��=��%��~ n��S�I@OGCh������a���H���܇�"xe�g�r߮���F���1-9�r(����z"F�v�����-(�O��_��3<��k���A�s:[����J��N�.�#���TC���o��f��b[C��/�_8u"�LX������	���L�w�+��;b�dzA�[�3W��W�س����	Vab��ԣ@B���SQ��jmoh����͚���vdnn�������I\�g����7"v]�\�W����r�X��yJ���c��҉I}����_ٚ�w_������Y��M�A�Q����#�u�|L�Y�"��w�!�9	������gLyO[�5&O:�T��?�Eq2J�d�5 �-ӯA������!82M3�}�L��/T����;6tpC���W����I-��6���)�Z?�O���e��9-7��7�<Jm�����eį~��g�O|EdJ)i�"�0ߖ�!bA1��=�=�ѫ|��*�V���/���8=�n����h��ՎI^�<�e��	����4w��^;Q+�Z�{=U?�9{�J@%�O��� �J]��<��|���8�KD/�%�*�)����
���~����!�ok���1��5���dJ�m+ˍz2�g��;!�8�p�jJˎ�G��1Ҿ^�e���
^$A"��ߛet�t��Ks�[��W��ľ�߁U?ZX���%޻�P�����&�/R��		�j�<Aݔ�����U鬌��y�{	#��I5pO^���Α,H\�٦̓�E\�v}��1�mF]�Y��>�$z]�ї��H����|*x"��/ ��X$��M�UZq�m�T�U���!�[� _d�r��\L�[�Ij-�g�3�Q*�a���FO
�1NP��x��I����"�8����@;����ZO+��{8�Q-�h>w�5?ɵspﱑp�:�c�����a�vW����3��%Nɩ��bP�r���GY�d)z����k�0�{C�3���.H8�Z@s�c$��&� =d��Wa4�/S9������r3D��N A��o��E��0��Dş��˹"���A�f��|8=�� ��w�c����u�=��.�dTz� =���F�J��x�����������1����hI���h;?�E)^��3�`Zr+��o�K����������s�-��^,��"��V���pa�;�'�W�jQ��g ]��$�8ܐ4� ��������OS�K�9��!R@B�r
j���"lt?�Fl���6FC� I��ȱG:�|��A�@S\,M*��Wp�W �����A�\#���4}0�UЈ	���������$z�N	���m�R:F�֬�gfZU�`(�Q'وF@��2��� ��d���|xq|��>r�u.�W���V35�����8Qb���<�g�V�z�r *�/�����hot�:���|h���hlx`/�6�U9y%p_3-��$e/�f�&s{�i]�b�� g����Q��Ng�~�2�fi0pa{;W��ɿ�iY����5J.��j�)7�n;TL�׵��!�è�J#�|��oL�9h�_�$�<9ƚ��|�#Ѻ��Ѐa�kb�}=~�-\۰��$S/��I��w�^�EjV�����!W��KH��E�Q���G<��al������A��5����"�YvG��AP�n���U1rm��zK#et���ڈb �ט��(�+�M�i�Ny��Օ+Q34�.i|#�aI�������f��n"|�5c������c�s���R~�iJ�慮B�D��x3��X�mć�а�I��{-� ������nl��v�������KױM��󆪚������)`�91v��zs��"�Y�"9v!3�7U��rU�Y��Y�������t��&�W��fN�Z�qi-�w|�p"�-�L�a����f'��B�}��2h��f�	�Ϻ�(�.XX�_968�Aɾ�zZeP%��^6]�ؠ�H���O>��4�O�T(o*]�����щ�]�)	a6��Cy��r��N/r�L�ԕ?���
�1��ׄ?e��Gx��0w.���a,��ruxKcͻd8@��W{ر:���4����Z��\�aq����!��eS̤Y����,p&��T�C	ö����ɷ_n������(�y\��̼��{YW��rZ7����	Q�s�`_��Z��i��z�+-��&��SiVS�(��\4� M:8U9r�J�L��Do�*8��nd�(��J3�#﹮=F��M<q��/i�d�����m��	e�(�[��H�
K��dII*��vl�-�!����.I��Yi��}a�_�&/��7�Ȯ���1hy�y�7�S����b��$|�*5>yp�`U1���J=��>��m̫�[��j����y�e��7�9H��PP��Ɋ�g� �v��t�Eнr��=���#��r�v(R�6F��\��mz�����Δo��[��p����\F��r�-��p�)�H�_�+�F��:�H��_��Y�Y�Q�"���s�-����_I�����q!] Phyk�+VKP�Ҙ:�o�����_HԲ��ٶ���h�����+����+Ϛ�ieB�m�j��xpp��1E�`2��vd��t��@�:�-���r�� s�@��Z�gJ;ϯ���ԣ!�i�8��þ\��ӑ�׻<�<�K�~?�gƯ�!��4���o��MX�D[C)�����"���d����LJjT6]�TJm�ި/�����W�������K�v�}M�[S��ck���Ÿ��챿�:9j�VpR���Dg@��f�6���J�q0(_]�����I����.�����C��6�-��!�疭mO,��x�BtԎ��fF\D�a����:��^�4�b%�6	UrQ�����?�4���R�I�ߙr�Je�-Kw�������R��9�e�\T��74�׶#J���<��%��M!9����j�O� ��o	ܻFB�P�m�I���Vɺdc	~}����4�ǡ�e����I<��<T�s"��S������!;f�ߏ�q��N����d�:Ʌ��ͯ�vK_�K�w�L8�'��u���y�u����&#P�a�N���%+%��J��T��Q��u�f�~ۑ9�tr���rG�xg�T�Ԧ=l�����(l�_� ����wMUI�ַ�pkW5��5��J�/���I�!��o����a����I��o�@+����~�_��2�^����Y��}3>�*�īQ��������?L�@}���)�>�#��,P������q�/P����� ����F�z�Ѯe7P�	�� �s	��[E��+Bz�V\�(��T�L�̚���g��^*�W!|ˑ��x�8��{�$�K����飃�`��hs5JC&�޳0�\1^�0�p�Ĩ������mB�/��اb�L�!�@�`8uG��%��HȮ�9gO��E������R+������}6��5<�c��Q�mC�$��-�}�o>���*��NSL���.�9�e��>*��A;)5��Vo���`U�>7��ld/���/S6��y�t� �IS����J�;����+��X�(�qB���{�jcn�D��7�3F}�������>��7��~N3ŎA��T�ˏ����iG�5z�+������BV/f?�.[�T{]N���l�N������{�V6�(�������[��VN��X���	K[�S[��c"Eڤ r?�cR�X���G����r�.T<���O�Y��H6d��`!R��g�!=MoJ!-vcc&p8�*�&���� !����n"�ӈ��y���؁�!��� nd.�}Q!����K��R\<��b��{��ĝ��W��y�@P�Iޚ.�K�Tykò������y�A����\�Ԇ*�i�	]�}�+�A�A��R��")|~�"��{K4�Sг#��;z�&O��po�i�������>������惾vԘ�֕����^ŵ^��J��PQVFC��ČF�]`�Fĵ�}Ó4���3�3@3�9F�gXT�2=�:"��F�8������<io	)�驎�+�B�|�g�6:�e�@�@(����6��h;o��̥���iq7-L)����$�iO�44$L;*&E��*̄5�@r�{�_V�wGl������Aˁ����w��	 n^}��=6�j'W�Mt ݿ~��>3�ʛoRњИ5�%��\�����0���Ċ������-�f%�C�&�}�3jBӡ��N^�e�5E��og&������'��(��<��)ʐ��2��K$�^o?g!��v��{��=>]n�?���pen�s���h\�:B���x���%���BU2��[�'[�3�3�ߓf/6�)������w���!����B�ė�/-�h�O��5�G��y<!n{�Ao��5#��^K]W� p)�`r��Ś<����,��\��Հ�(C l_&D�5�0�e%��%S�B�'�RT�����;yP��Щy �ç�)�	B�N���$��1@&��ٍ>ϫ7�-���Q`�B�"\X����^����&����� ��{��a��AdTE;��┟��6u!����hQ��+��W{QͿ��+�_#�ǗA�g1`�۔�M��X��<��RJsk��cߔ
����56��B_�[�щ��D�%�x�Q��� kŗHs��^�6�䔔�&�#�(��.������&��V����m/]���_Qp�5��*d������sZ�����oSb<I���s3�Ո�'�b�'�B�,]6S���h�G9�b��:{8�*4Q�3�����K˯�p8�Oa��JtB1�7�mt��VU���h8��K�����VuG`��g��Y��Jm�R���o�M��GYP�8	�.ߪ���I��d�^�ƯBݿ�d��J�Ygd:�$l�m�J�H��s�+=:MI� U��)l�GZ��kc�ŵw��oT�zB@^��
._{ȉ��b���Z����ɸ"�-��@O��e\2�E��s��`X�ϳ��bZ��M-�/�LZ�S�4�q�z�=;��b0ł!oZ#6��@t��wM8٧�4�ڛ��[���F����Დ�1�ܿ7�����G]���b����(H��B�I��KM�,��t�1m�,�w�o*3�Z���x�>�����6�����T*��~�N5z�YB��"��� O2����@3�鯿v,,5��2��
ZJ�Z.�
�K1�<^�
�m2S'Z�j��#.T����(f�U��(�����S�1��u08~����_�!�z�=��X����#]+��+���O�n�m+4\gI�Վ��ǪT�u�i���R�29�h�bx��r�S6���ߣ~ ��e�,UYܝ2��t1���<2޷�󜅱�-������"RՏ�����Lu);�G��P���R<�.�V�9�'�ϑ}��е��ƨR'���"�l���{|ý�A��I��`/J������/�^l$��֡Q�m�f���:�{�t�lG;��6�$-�����p芀�;��'����~NkI�V�8ȥ��;⟒�S�I�p�#���ȩT�I"�n�j{�ԭ��x!I���{���	�!�@�MlLZo�չ'G���R���6A�[ۤ�>�ᬔY�#g�e\J�ͳx��P���hWH@ϴ�Y"�YZZ��T����,s�+��F�1M4A��r�� �^�[��fH娑��h��
 ���;�����>�w[�+.
�~�Daa\�[!V��\؂�n�$z�0�k���'��c�s�^He�AN��~�u��m�E����R(m{���粦\S�ډ�KI�O�m�y.A-�hȝc?������jg�ï��GT�O�V�5�kl��ӏ;�Ӥ$��u���w��m���G����_��,_6g�3�+O� ��@"I}�O�3�{���[}} �Rkm���⚞�'��lW�nD{Ɣ���� ���ے}����H����Ze��Ԫ�z�*��1DH���'0���8a�E��� �q
���s}n�kj\8"Nm����q�K�TH�
�Q���-�����uCFF��@/�<+���s���k!f@�lY�i�}���I��ؿ��C4a�Z���FW�;�h:{%��|�U/�&
P=Z3�Q�Ԫl�lt8H�����ư������&�����iQ������� ��r؁=�~M�A�t�bk��	ܳ�S(H^�,ʩ��;½��IxR��<�$�>��$���[=	���)J��W`X��7^:��Y�W���nn=F��X�V>����\�/k������v\���R�(�4Q{��ӈ���c={t�?P�/^��Nā(���묮� ��~N�{ɉ$�M��E�b�`��3ش6�cP� Hǎ�P71�"�w�������Ê��3(j�l!ӛ'��X7�o����:;�;T�h�\�*���4�P�(�:Yk��HHFwD�!ڤ5���/�>RzH��bf��Kq����6�)Ά �b �G-��Yl24ݷU��AD�o�g��{�e�<{3T;Y����`����O#����>�`�fJM�p'��hѢ�{٬���Z1�=X�u��˔����L U��0{*�J��rt�s����'::����g@j�uŕ�hG"IT��ўD$P���}�Jt�c�,��E�J�-�E��ɇ�_��~p9�ko�;Z�o%(�]�@�KGbE	�ʭ�VjR�bu�m�J��%�ǞCg��(�^�
�;�چ0��y�Sf����;<�6��*�B�y7�����M�n%��u..y�.�u�\�]��X����=�S_��D�ܢ{yv�w�=z�,$$饅���(��k�[�p3�p��2�Söd�i�%iKP�����Y��Z���y�45p��+�t���H�f�u,�qꖜ�z���H���� S���Y�'k�C��g�y{��Kk�e����і��Q�߻$+��A�K�0�K{;�)��&��6yt���L��K�,� �����=#�``EMUTr��=��P��Gk�[B����whԮ���?�<���d6k��G�0����ب=�I��,u�fиBf�4d�r�EHW���@�Ս�{�/��j�k�᛹2@B]����4J�*��Wq�V�SR�e}%귭
�U�ٜj��}毬��D /(�H�[M�N�]��H��P"����i)�S�D�W�m~N�^xƹ��L� �6���9�M	��8^�6���hD��]n�y��x�P�ĳ<���b���:���z�G�v�2�T�n��sa��T��Fǀ��)s��U<F���&J�8��zwB��~@���cca��7�h�E쑻��:��|�hl�b����:ք�j/���X�\A��ܪ|�������e��Ms�=2.�6L^N����3I쏭�qI�erv�U��i5���$��T�v��]�GVq�Nm&�Gݙr��g7��AmYv�^+�`
X�%@B�����/�i��K�@gm`�b�1IPN诜�TɌGx�EˁW�|��C����'�捨�����c����Kg��*Ϊl_�K6v9�˂gв�Q|e�\�6r���./��|�Q]�ݾ֐+`�o��"@�ò�Q9UW�#VE�"�'W��� �H�d�ұ���9l���=Y��8a@��إ���l��v&��J��n��X���ri?�k��CAA󽼵��*�#
�	�ܺ��#�	��\�dqdjṍ��� �q/,ѹ���ݢe���`�^Ga�o�`}��Yt��� p�����q�o��p�̻���ޒ������4
�Ǚ��xb��,��3�940�S���6{��=�����%�B��^U�T`dDGysFX�m��
�A��T��ꢫ�0�}���~�%o�ǵ�$E	w�~2t"��p�V�O�Q�N�TO�g}+4{q�|�����1��0-��4�^d޵&E���+Dr%-S�+��f|�4s�hlML�g�=�Sq�4���X�J��6s�t\����PJqC�#	8w�FF�Ӌ���:B�̕4���(2­qdL�毼�6��[��-W��iO�m2֊�aƒn�ww�ȝh�yا�l?&��e.�/��h�7��i	�$�sWS@�*���5��+��D̞6���S
P��]��m��s�^��ׁ���tP�j:����ƣut��0���;K-n���:�ru�>S�=`�Y#&�g�B���Vo���F���h��2|�p�������	*��.t���M�w��3|�}��5P�J���a7��܊����<� 8��OE��[�"-��I���SLu@����fζ�E���w�e@,J ������	���ˉ{�<Q�$�j�X��褚���E|iı1�����
b7uLxt|�F�������������� ����/�rE��=Yx8��$<����Ȣ�6��̘n���a�^:�A�z�0i�!�Z�ZG�[Q�V�F�H�)G|����u��'���	6ڋKd�e����$�W���{VC������Fj~��`8`LT�������ӣ{8��Yy�1Yi|��;I�c��QĨKw�ý��
����e�����f�tApk�u��Fy_G�!g*������G`M�u�i�6/<!�=��f4M�J�m�����sf�h v���d�QIiz�0\H���y�F'u�
h}����7s��,�|U<��j��fU&�lp��uѣ�a�G�g��z��2��ƮzM����f
)�/DCZ����P@�1(���\
�,�=Y�N��P.�k£}(�<�PX�6�����n�����'G�F�rX4)��ʰ,o����ۑC�=����KV�#�%6��32�l@پ��5�֛�	�鋎�����.��p�����R����-3��g�Ǿ��P���q4�O�9R=�ї굼^�o��H�-�{�uΣt9\�ቌ	͐�	Z S���D��Nxޜ}�̂ava�+N�E�ۏP�@g�&0JT��s<4� ۙ����c1�e�1�,��!y\E��l��CH�6�SJ��(��Y�{�՜f*���*bZ$:"m-��=���~����lM@-�/�y��
D."|S���l
8@�s*8�q�a���)d�,j����3�ٿq�E�z�k`�Ű܀���Sn�)�M @f3h��z�����K�/a]E�_��M������%z��2��p26T�W]��V���G���#	�by^	�����@��C��e�w�C����N���6�/GN�f��0��)*����6y�b����x��R�[��лS�o5�|El�
��������8��_�<���������A���l�-�E�QJ'CF�Gɷ�4�=Z��9�^qx ���*�jD�Rc����vGeR��E���@�,�5�m��.���˟�ݦM��EJ�Ԉ��V�Z\��&֍�"��8���t���8ͭ���%��K}���$0 d��΃~�`�M	��6�_�����c�P=?�)j��w)P���qp�gS@����[�_&K��|���y�R�Be�}#�X�9�9����L)`��_�������4�Fϝ~s�
���hSfT�v�a�X�]us���)pj(�xA�!�"x���3�M�C��3&��옢���^.6�]�6�΂���P<�9㫩A�Ŝ�C&�\�5ZPie=�O�\��� �q��l��:{~.��3V-���^����G���ގ�F���}17�`�Ў��"�o�ͳ!.�����>����>�L��Bo�Eԇ����qI Ӡ����H5���D)*'����P���E�ɦ����#�	��O%�'p��iʦ��Ƅt��b��|3�9ll���Xz�^���j�ؤ1&���_T�5cՒI�μ�s��)�g�}M^���~��4B��y��ǹ��T����;�N�Z�o�L.����C6�B �2�"P���w@�a��T~��OË|d&�_�` k�j\�ߒ�g�v�2w����B��/f�Ld��?���;���WiL���4���s�����M�Nq0��	a�1���~�?�
��� *V�����FM3.H�*؝�� �bW��y
oW�� <E���n�#������gSzR$o J�#o%�;�H�Ay� Y��2G���󳺍��x�v���T&	zL�k���~鍭�p愽v�\��DCz����֝��O�<�o5�~[ԇ�����4݁I�M�ݑ8�H&{*p�G�k�F⵳%�JT�������6���uХB�f�x���t��;�J�#���@�G\z�?��BW����������>�6�������O���~R#��2�IE�Oe���A�M�7���FA��
�Hz½�Ͱ�>w!v�{��;�_(�c�qzF���k���n��+�ҧ�W��5`�%8����a�J�CU�������Wp�P�*I�����ʻ�1�������\�8반(!�T�)��r�;{��&�h~�O� �ū|�l.��ڣ8���yb��[\�u2`綫�'8[<� Y��Z����Z�K�C���@��*WL�&q��|�o5�I��Y[{O�f��2�q2Wb�)k�qxjJ�/��{&~KtI-���wL�@XK	�%}st,� �? �b�Z_��q���ws� F�����]�6\�y	�I�J%��Gb7��7���n|l�͎�%������l��XI�{ͼf�i�.�@^�ÉYU�d������U9�P]\ڥ1��T?f���
	��V)b�hZ��5.���ϩ,��H�C]Aш]?�XU�ܹ�i϶�~��0�
ֺ���YҪ~wc� �B�2�qV��C�+��׍�C�q�:�O�į�ҎN�l
��D'�e.���ȋ���) ��y���:|&���м�����-Q2���,EL1���0�=~���P��p���!DC�pQ��bMD�W�t���>��ɀ�AB��7�c=�=�~���P��<��J`\a�j��V�	�{Q=����������ʰ��W��=�F��8H�{SL�}��7��a.��(I��@$��Š/� ֡�����ߧ��v|���-'�*D����T����8hφgDp��l<|��HHF�I�����5��,k�/�~9Q�L.����$�W�x�!+( �9���&�|v����{�:�}K	�R�9���;wt����M[T?����RW,C�IMx|s�+�[K��7j���E�lw �F�'�Ұ�$�@�c���+�?<�&2�}�q��g�Q�B���[�
x!D攅!��ֺi�o�J⾇�}��KP�E
����r�p�p�	E�\����\`�[L��D�O��B��	|ْ���/�z�2&:�i!@A��CJ��ǗƑ��c����s��^����;U���S���A��&�����Gш��"Ih R� �{���6#B��0�	Р�dWEl��n�����ؔv�Wx�x[�Ա�F8>��ʾ�Z����U��3~����`Y�?�� ���H�u�Fs;eW��q�-�8~� �ψ�;��"�����SKj�V�%E[8{��fqA�d��GY��@.�j[�[�}ur���ׯ ����$&�U'���%�0���XqǑ0�ε2��Nklp��b��R1w4�V�|i 6
J45�^�wMi"�C@D&���1۷�/��P��U�pcU�V}3�̽l��1l���e@l�iqo�D��Y���`D�܂�4E۽Y�9֒���H~S�hn�}�T))�5�!f���f��(s��?�}�>
�B�m�$����������YX&/2ܞ*�L�:L�L�s�Y��J'��Z&J#x���Qs���|���9[H��QBm]8��4էT*dW��/Ľ���i4��))H?t��p"���}�!������\�Θ��g=o��a4u��̅P8�����ޯ�������[���Zh�c
!Nw:���
f����x�ȑ�-��������{m����"_�	Ă���:�{�Z҄&`��V��:�U��#垿Qo��i�VS-���WJT����0��ϟ �>�J���<���%��+/q�7�E�ܬ�H��rZ�M��s�R�qCB�WA	j���k�[�'Y�a}C��E&,�9��S��e��#��$�)�9�I0��K�i����w�)��E|¬���#�NrZʊ@aЍ�}Ҡ��I#е�3���������k�ܚՀ�8��+��� �F��>�	L�%$	�ø���ZϢ_k�ޠIU���BW{c��/��Q&�D�ѯ� �&�`A�U���J�2Pta�ġ��O����7�/�t$9Z$9P;��r��R_�#����t��ݳ ��t�|�Ä́-EA�����T�e�����)1��a�����[Ap�>��@�pk��h�c9t10�ç�+Dx�w���9]�%>�ۯ��E�%���4��G��m!���2�����c��t����e,�`z��K'1E�v0ɁJ�el��v�m|9��f"�Uw1�nt����zF�f4�YĘU�4t�[MZ���&a&��{�!ɏ:p��4(�U9��a�Hpz��u� �tt�a�cL#��2�1�a�!}�T.��_9�2BВ�����;$��6�|�3���������rK(��~@�V�+at'q�%l��`l��J��'6"/�,f�y΄˿���I�w8�1Ǭ��e���)c!4���f��&��C\S�=.;���R�~t�kB�c����cr��"�`*��??�)���6������&�<%��D���Q��p+e�2�q$����'��X���� J$4�ȼ��������,��^�<��l��&�.{;����Ի$󪚷�i�֨н�D!{i.����'���2Ա�H��8r�uz:QE���eeyK���k��W��g����.tiU���GPp���$��<�Qi��p|�9�B�D΁.�j�s.5O�'��A�;j���W�+]��gyl�?��ql �@�y~�G�h��h�Z)V[���͐�!Ҩ9��oO�@�yP���xGu[Q��P��K��[b�L����ڪ�13Y�D��^ã���hI�h�X����"=���҄�$��,���}BU]Xa`�����$�@���߻'��pg>��rq08́"�lY �`�,�,z;�|��0��"�*;g۝|���g�p��;/�c�ݒ��v���˪�����Z}�K���$��n��D�:�RN�[�R^(�㭹K�G�Å��>"+�G������\2��H�l������g�%��G$)A�m
NR��Lx��������mV^��1��FH5}}O��q���o��j����5���/"�O$�f_g�����XT��M��wvȭ_|"�ZH���<X�)7����'��m+MZ�Hm��5L�H.[({Q�W����9��;�;,Y��֙_V�����M�6jN��嵚�m���yW�m��E��{3��m�K��~늂��R���2����*���0\�����+������-���`
��̹Qc*�B���^kb
�W'�k�0���r���Ɍ������2��r����ފ�o�K��h���>V3�z��H�,P%�� $��8|�Q���u\�	�j%�g#�ɘ��A����d��J�#!���Z�]l�oV�\��/����.�&�"���9��FW���'}���f��$�,B�i	���ը�]��U,�'����A�������G凐z�>��W�+��5��e�����
���<T�J��
�+Q�}��� �G�Z��u|�q�8�L��/ �~�dɀ����c۞�rh�K;#�Y�B#��<�H�*Ķ��s�i�|�
X�����w	h���`-YD�w׵���̤�X�aF03��<8�z�h����+Ae�ġ�C��,e�`��NV�R�Eٜr~+2�/B�]9@�SP	�;�o�%��K�n��{��%�d("�!cƅ4���(6g���I㴙 .��Z����4�Z ܚ*�Y��h�o`���`����fPAb�W��Bt�3�!y����x���ۂ��>
������$'�g��<2 ��l���r��[ N�k�mh�L��d��gK��mʻpP���������V��b��1�b2�M����Ӕ��ܙՑ��Q�O��� P����6�R�͌�;u���=P,�Y=D\\�8�E�@��[Wv�o��2������YP,9�/��ԙֹ��d��(���ޣ�r���,Ͼ�0����҂{���QPg���3.���������굦��7c!���I��F���$�L��t7~���8B+��"
�e����Y�]Wj�2{���Y�S�O�%`y�!�A����8h2	�j�t��
3���h!�+P漶�w���>���,�gߋ��=����G;�n����+^L8�/?�"��y��[2��J�G��a�;n#��g���M�;ئ��M۳z���[�^|���r�^�b�W��F#w��M9��׬EP�}mm03���QϤ884�7�ߗ+��th���z�{8R�JL��	Ֆ��䦢�[�I߻}��+��J�G��S~�}	�V/O�_Z���M�;	4AO�
���߸�
��1���1�����n<�l�H�'�Ň��Ȣ��`�BXY�T�t�D�
/ �:Te9{�Ǚ�['�-��(f�p�E�#���1!4�s�,˺a�T�=Zt��o-�"p�����P���]b;� �n(sm������>�M/qS���O\c�����ĸ�|P�������}��;e|�].h���ߟVƛ�ګ$4W[M��c�x~�*r��m�S�b���2*�޴ ./��k�i	�$ZT����R̃,���)���굫�0P:&�+�?� �K�,��
>t`mJ�S
J�7%�����)��
�H����s��� �a� ��y�wFlM���FcGRl��6��B�=���?���M���WЅ�!3��'i���m�	�B�%��������]1ԷfC��y#���/����g��ӧ�@�.vS{i��K���:_�1�L�+�QƁǝ�;���ȿW��P�*��ϓ-.��8����!�n�t,��p��Ӹ/�3~!����Ɏ:���I}��������I6�("D�̀�[�웢�>21Du�sdƥ�b ���<��։���d��S�5S�xj>`�'�S���e&5��pfN��O���B�y���>�������!(���������C	}��>n��Ժ9���%U����h_��c�XmW{^�~��#�j���#Wx��ͦ��/��j�|/G�F��_�JM����X7�P��o8+n�p�gG������'?��+�[/#B��VE�=�[�f[�=���@m_{>
j�vd�T}����Μ��k�m�'��@�^Ձݹ���bah��7�����q��p��>���@^q�����'Ơe,�#�؊����(x5�.���-�G8
Ι�U�N�Q{V*�QD")���wu��#�75���Fk���l�,E���sL����rr��F_�8�� W7nKn�p{��91��"�f�Du��'��RFp� �y��>��eY4�ťEq�YzuX��e�#�_�,�ڰ��/t��(b���0	���ZI�ǭC���THٞ �mGyy�ޟ�K���$V��������QyY�*\&�J�����ҟ�|��/֦@Yr0�*;ض�Bk>�a�v�y奜Zl�C����s��7�-K=ȍȂ���� x2gw�L�x���SQkB��u��_f�5.F"%	�^� ����yk���꣭ nLj�2��l����7�
	O�6��f���,�V��yj�(���Ab{���$�^�Xsb΀��=τ���R����9���S[%��!i��JC��mƗ�:3�і��'�å��^J�~¾̻X����H�ۜ*��!1������gCn|y&u������a�D8��?\Zff��3˿E���=�ōG9k�sr�y5[�0Һ~WЕv[��h�	1Nnߛ��z����@41*Hi"&�S�N�� ɉ$��s�P2E���������T?%�\��iuC.��v��-��#6'�)O[��K����joN���p�q('.���p�t�Ex�Y �:�'��}��j��̜j�vS���J��'(~�*[=�VJ�5�m�}��|�p*+��.
��ʸ����c���ai����YW3�)$k�|Z(�9�llZ2�;�D�y�n<4{�2QiRƺP���gp�� ���Ԫ����4|.�S�t���o�P�<SUy��}��If�KA�5*R��3)�S'C��������_����1
��;Y�?%����n����f����f����E��3$/wo_�DR�Y�Z�˸B+M�|:��!Ɍ�gH`��`)�N2ȯ�z����GʫNR	�876�H6W���ω��%6����m3�L���v�B��3�m:��FDˁ�(�+ūM����iH�������6#�-��5�j�ϖ+~q��a���ug��P-[V"45S��X�nJPqf�I�1Z�<��M�k��������b���}�jw�?US�;�+����;��Nuu��S8Y�����C
�3`߫���� BV����tk_��t �UN[ϔ�KrhSn�k}Y~ګw ��;aF����c$��{Z�;K��G��A-���"p:�x����;G
����z��u���ڻd�Fm���)j0o(�7��������]tE�YDM��u�El=�	IU{1��Ӯ����
����-j�]$C�h��l�.�ڞMYu�@����"�C^Tx���O+>w~�j�4��܊Y���X�~����`y[O�
�2 �r]=���.�s]6��pڀ��Gm.�#o��C�Y�:���*����r�]�JȰ/}��MB�tP�L����bֱ1�LB_����t߳�^��o�l��9����_S]+�J`+�����<xWʹ)x6n� :��k�"�\��v'�_;����j�����a5�*���w̡@�нeT���fLYI���ʦ[�뜲H�a\�a����[
l�ذ�#��.C<
����I}0��0�����O��7wg;��MȽ#����4�D���x�k��s>�ʯ��Am 
���>z���W�z��}�V�t$���"NA��4�h��S�䁼�a���W����C��&wg�as�.G�g�럃�N�ɹ�m�y+̍J�I�f8���ê}B�|v��X3O(�ع��%s�Q�쁑ήC��M���&�ν����@����cp�5@�{(�[Y1N=�|�WP��O{�z�+�/prQ�e+�Y 
=�&/Y^�-w�'�0V��>g:�A���`��v��#�aW�FK�0���񗵬��I�D��g_�Tg�C���B(�p��H����w}������yq�X�:�U��Ł��d2[P���LDQ�(̀����� YY< �Ԩ�gP�y���O�k2�[Љ�\48���x*FSR�gc�O�n�ud
���
����J��8wc�',���&7�O:���oG���2ĉ�0�X?���^��؝	��?��J�g��:WE"���_p�y����O�:�+���,���||�)X����Qtg�iBQ��>�p��Y5���Y:��+Gx1���8J�գ1�o����}j"eGu�R�S�R��,4��PӋh��ӍE��H��,W1~�N�u���4�Sl�P*Q��w'���=�
�3 D;�k��6�:|:�X��V�p��� )�vE%`��d��N�P�ޜ4|�oS)}v���S�I��QfG�m0r�l��)�����-�ﶤހ��_�Ƴe��#�