��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� �4�Y?�5:���팑�����=��pv��ξ���������l����5�����"�|Q}��Ω	(-�c���|K�����>�EK���C��R)��P�j$���j{�*S����l���M�P�e��m�iA3�B,_ @���@�}W��"�.������)Eձ�=����ݽW�=��|��3l�VL��$�ءf8���xY@²�/DK@���s
���\9g>�\��ir��p/��O��L��"w��}sR��wt��Vh�I��V������tb�Ѝ�J��,?~�	�lj���ӆ�TY:|�0����kcW��H�y1=(��# Ą��)q�U%6�8�x~�qZ+s�d.�x��I}�mI銛�1�N�3�pKìb�	�x&��o��0D�;X���
<�Y�3��m���r�:����(��1��H���`E������c{Ё�I/y��Dj~�Ķ.�T;1��F����ǝ)�CˍPN_ߖ6)�����Z[�?s53f�0D�ϟ �߼��΄kx���W,��-��M4F�[�����Oa	<�R��:��A����\��Ƶm8�b��$f���QTC�X�@Y�=�՗��W�1��_��"?�{8f�p�u�q�#$�pD ��u`4�Z��k$(@����_¥�=�R�-��1�R�ە�ޠ�2o�L��B,M�Ih��Pe�LR��{3���F�ʡ�������j�~y���OY��gE��}�JD�V7���!D�ɁJ.>Ο[T�B���UM#(c���w�����`����>ub,[�\B�p֙�b!�n�&5	ʦ_�W�)���fH6{$�I��#��+�F���P��SJ���.��U"(�?� r�jD`2Bп�C�s��cs�Tv|�p?,Nƚ�wx�X��;#;�K}�]� H��H��r�p_�3�}��hW{m��c�@	��8&���  j	���N3��B�,�)�� �KK%8y��+`�[S��66f}q���@�{�J�}���D(8�0ok ���=�'Q�j�$���� ��'gO{Ƚ�êE/�տ����d�J�Ĥ������?���w��)�X��A��i!�g��4D�΂�#R�椥@ĵ�h�n8����h��}�~������p3⠂�3WuֱI�����9���v�*��ʞ4_`G�� dp�v��8����3�>��?��z����ZB<l����L=�E�8�<y������8dU)(��V�k1٢H�1~Zg��811�#�}��s��t#�i�I,�&�M�+�gR�uJ��g���fq��<�*mF7�<��.-h��mFg f��B�8m�'å���\�cf"�F��@�V}�/G��m�y��)����3s��*.p�<�Z�'���$d���.^ER04�{Q�m���W�Q^KA��L*��3�$� qM�g~S�}��OE75oF�i]]�68����-��?x�䯝�͏�7���;��J��kx��9�Ϭ���\B�dG=��$�T��l�%K���W5�k�qx�����At�-��/������FnB�Nz�,�i��4^\~��gAcx�Ȳ8r�z����w���W�nU_H�B0w��*C�S	4Z��^�X���|��oG=��y�������֯����j�u��)of�t��U���d��aE{��Ɲ�� ����W�S�6��(��^��[��x�뺝&X	Τ� I�R�A1�[QM��)�񹒒D.�[a�3�67�Ug����7<Y���r�z�`g�j�ߴ���ȧ��jd�Ԑ3�h�?,w=���ϧ�`-F��$�r"������KW�y#�#�ami��o�Sg��H\�*p|�������������'�T_�Bj�i��#��h��JD3G����z��Q�B�w?HϠ����a/@H�Wb�}L��wJ]E�9���>�48�t�m��Q�(U	P?G-.�ˉ��"�����S��V���������j�nU�Q�'s��0N�n�%������V�4������1݉�A	P;�JR�ߴ��m%�� y?x"�+T/̲�w��ւք��#^f)1�����ܶӏ*?�ta��*C�xj�ݰ<�V�K8�/��tT�B����u���A~胏bT��0?/�f�Bg&� R�X��W�ʏ���p1�{�&S/�LN�mST�g����Es���S眺8�%��L��m�ejbef���9A���� r�j�^7�Q���q��$hc�>���O�8����V0BmS̳Y�ӎה�� e4�<��U�w�Y3T���*Q��Zt�U7:#:�[�I���U\�q��B�+��5*n-Q�f�/]8��
�����;���q�h)�TMH!<�f�~�?(�`�f�0��֟g���:�t�����E���� �[�7i@&���w.�UL�Ve�����L�������~�x��	�e�kw�(}�QDG�gͭ�q=�W	� R�YVx���J.6���[j�xs���f� Y�r���M����*龃V��%QxcA��]�UJ�v��:)��߂p�|M�|۽�{Z�df�b�I��+����
�d�[H\�a^�b���ᝩz�=���̮ڊ�l�uF��|�=8�nB9e�8T.���Y��^t\���l d��1�������x��l$����@�V7�Dx��z!��o{��b���e%ב��5oI���ת����s�h`0�ɂ���h�q�K�<�^�b}�a�E[�px�����S�>��#(�M�Z:�_Jr���S;D���S_r�