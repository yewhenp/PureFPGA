��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m��k?��V��6��"�"?�=�h�0��Q$V�=1zr>�:�\l���6�t���Qr���?�{�U ���D6��DJf�*	�	�خ����0ZI�=��?AN�?�{��w̬0�%����ˢJ "e\�5��=sڗ���h����6�<.����R��ł��t����s����a~����Ғ��G�'��������p
��QÕ�H�[򫏋=6?� M�=p�6sٞ�����V5fZ�1�ű���b_� Ҹ��������D?�3�N4/	Q��O�k0��<�cW'��k��"~S;�>%���[��S�>�d7���gG~�;���an�]���(�"!��tlA�"Ƥ�K���͌�I*��7,�N�hg8�3��:(�(�;����2YϟN⤯ER��,�j�
�&w<��y�w4"�s��y�L$;�ju�h�Q)��+���t\y��P���q��:K��<f�:r�ƙ?6��[��ڱ��]��+��:�����2	a�e�~b@�nm��h�	���\X&zX[f;�נE)L���Y7�l�'KU��)�%���0+�| �Ѕ3��3 ��p���3ȕOW�n�`��?Q��t!�^)9�q{P�Ks�: ����
�n2���2?��5�Y&p��x�Y���$U��K���G�Ǐ�}3E �W4S��e�f�ܒA���'�M�D�,�{֛�;U����X��c�WHߓπ9��֮1³�݃�nj7E�e�LM|