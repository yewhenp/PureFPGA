��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� �4�Y?�u���/1C����4�y�{�`�SR����@;l	�蹑�6#�B?W!Iu[$ZrK/2&q^u�Y��	�KN������K-���h�2��Pl��]�[?�4��.4D�wٟ���g�[]�@aGq4�հ�����9ORcmd�i��_���:+�]�t�b���_5z+�Y�m��$׳$R!���3����M�@SX@�a
��T��ZXP�$��x��CI&�*��3_v<��d♂��:9�w2l�~k]�������?:@M^�������-�����.��U��"끰il|��a�ŕ�8U����K��3�&f��8�Gڲ�9t� �ez^'ˊr4X4���d*���pM�*�2��� �m�	T=���{EsP��!�i�a+o���g�V/伅������^�Y2�r�\ki���sA&h
rh(��0���o��Tq�����h����>������[N��s8�1�}r��0o!�!IV)�G��	��4��^ou?�Vs���R��v����dۅ���A�C+<�"��L����G;�m�!
H��+:��Bފ=o�=�K�v|0 L���|e��Y4����%��Z��X�u��{���Ut="�!vbgB�%�ɷ߉+�'�����_::>�����������W�~�bC���g0�]6����Z%ņ�Aly��]��$�Z�j^�����}SUFb�t�U��J�����v_�)���M�`�x�졊����k̟��/@��t����*5�(:4��n�(�,:�$?�����6�{�����M�7[x�oڑ�-ꥋ%�˙.�}n� �ys�)F�_�͌lQ=��R�D�ˌ:n�R�� �ם�/Z*�0:er���D�)�$:�J�3*�/���j��.f��+�}�'����0ϼ����Ԃq|5��{ͽ���i7i\'�pXp=��'Ri�H�_���Z
?M���E_�3��6����3�:�X���>�'y��׉:XmXwz�sx�)���n巅ޗ.��6���us������@��� �\Q�Y;�r���@fazbu����߆&��[��e쪼�;Z�{g������%@]��G��*##�i0T5Q� �'G�v�Mdތ��:QF���������\:�@<a/ƽQ��9�;��D�<g�����\ʐuM�A�IxG ���T4V�˙tKcw1�H�B)��<�o2��c�sA`fP@A��E��ϰRJ�xE�ˑ( ��6��l�V,u��@��>�
F`>	;R�ԋ�nྗ���vӲ�t���8��E`�����/�h=���+__�dmja<0y&yl�Fi1� ��8"�L���B>���
EV>h( ,6ܹ��Kw���]:���z�E�5�T�Q��]GA<ߞȿ�k+,�䜫�!�ߤ=Dӗ*�4p�M�첵@k,6{�����8��>8�8���-:fz�7������R^-�f�XZp�{H+���D��MlR5�(�)��{D�6D�~�U/���+{���U�.�Q{�$\�:�cq�% o^IZ��5���R�@�YY�h�=�Y�oxk^�S95"0jm����Qfm��%;����'���'����y�庚�S3�^ܠ�����[��((]�� ���i,��h��0콢ݵ'���z!o����s�ջG���锈q1�䍾�� +���XG�R�|�9��	"�I{9�� �L��z@ʛ�����#u��!Sv�pW�K�M,n��c�&������ɨ �Ƅ�h��,����&?���K-��UD���}!j�����^�nOؓ���4�`a��p1�΁_C�ưd����(օܚ�ؗ��Z��/�k�#WR-�h$u("�H�'[��/�]�w�;^��{:��������?�<�(��;Ac��U�4�.�1������d=�=f�.�b�!��ƌ�+��7\韙���ޓQ�%�Ӫ�]��j���(�Ɖ�Zj�|v�Yz����\����5}�( Z5ǳ������OTD����S/%ӦQH��=.g0�3E/{��x�V�tv2Z���`R����H��>5�����q-�?@��;���oCXn���p�Q�