��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� fg������%3�#�����-4/�__�<1y�쮰�W{"	��Ȯu�Uyif&��}4o�j�4lLl�yʚ��Z��*��;Z�z��5x���t�XEY�S�LԋU���D��7T�$pL<~Yt*Q@���@Ӹ�����V5Гm���)�7nx�ƭ}TF ��MJ�Sܧ\Š��\�;�.6M{��8^��N�*d\
�@�a���4�ˀH����ہ��x�&v����]���^���jɘ�N������N`��l��D���z >˧'�A[�l|�ר�N���r�B�_z
L���&�Å�.7��v�5��,�l�ѣ�a ���לR�UɈ�.����d�=�\����A����}����,�����;=�)m0vfU�9��V�I7:�V�F�9310��=F[D�+��^�����Vo��(���P�/�^���v�ˏ���k%��[���7W�J��6n#�;_#��3s��/���c�_%̧l���91U��_@�J�T�(���0`��ev���LD/�+�Nx�B[��^=EV�u1#'�Lu�O���mUO3�����s�U����|!c�M�R_��s[����y�`�Q���>����dT�.������JO��������g�?�j����%����k��ؗH�T�C9;/?emVN�|/�El����h�R-�<t��L�)���r������7��A���@�-�k���5'r��?�l���v�6���c��/�W$���6-�l�ρw�W�o��s�+����Ҳ5Q�s���'�Or8F��F��Ӻf[z{���ηgj���R���8O}��Z�T�?�D��Sb:�}��$ȯ%n,���;���;�gpE�e��o���;�%��S<6���w	��D��z��i�Z���x
�/��Kus��iv,/HGO�%-4�$<���Ix�٠6�ni�_� ���b�Bt�����̬3����%�z�霰����z8���o�ӹ��`p��wͷA�wz��Y��+ݥ�R0�a*�_Ԃ�����\ll�魉� 3����/�|��opb$W�MH���M�_Κ�j�:²b�j�S7t�'���ޟy]M����}�V��` mEܡr�a��>?���q�,����E5��jR����F����wFop=�J�*S�-(���Ә8��#j$o˄=�}�ubo�kH@`"]��z�c
�O�[)�;v� XGha|t����3O0������&DNN�+�,���[U�Mk�]y�kE�nJ3"	�;1�P/�8��p��A��`F�w�v�Kqb~tQ`ǹ�LM%v�)ޑ���b^��I�{w�69�x���Kъ�jhĭ�圕�b0i2��t,ߏ�������W�������S'^�z!=a���B���5��c��	��,�~َ5���xǾ�/�$-��ajjw��5)L��ƽ�˴�5:c�Z���V�)��1i����[*�x���;���2��	kˇ�b�1���������kI�E_=U7l�sn;�Z)	v�����;������m&��F�V(�g�Z�g`H��g�Φ�9$O��J�K4��7,g����ɕ�i�����J��?f�?wbƏ�C��Z���UWq�	ߤ����e-e\Ň!��㢳 �2�ݻ�C��5�$"�c��Qy��^�������`�x����U�'NJ�{t�Ykh��$�8�&q��l���4Hj�:��A�!-C?���mdzG��-(V���Gj^�x�L�&PB0��:���H��f�����CbfCW��!���7W�"�dZ���亚�E��h)�Hj�8B�T���(���f}��X��,$q�f�b<4}�@�ɾ���{t��lL�b�z�a�D�٥{�
b��I3�����e_�3d������y��(�:3ٓܺ��^-6��I��i�̑c�!���WQYh4��Cmz�L�M�G�bT�j3�M7�����Y�g��J�?��29��>O�6-���8}-��i0�rs����I�ypi�r��G�[�9gC~�spq	� �E&7F%�bv*Y-=l{���TK|P��E�����*�@B��JH��s<����$�#�%6K�2$+{<�7S�E��^�tO�@�H���;*T���7}�L���Ŧc0�dvA�1���'��"摞ʘT��A�y�4p���U�3+�i��쨛_���%�>�.�[m��%d�o/�Q��g��Wy�F��/���%�b�8yL>�?r�N <�eف��~'�HX�m�9,`��x�������Ӡ�y�*�}c3�D��ؽ�4<�98ye)��]�����3o O`���$�ȷ����[]$?��Nw8@�b��mv� �o�S_�V�^q�!����G7�ּ��}jw���˹`��?���e�L�'tf�]]%	?�	��;�R��ˢ�_:�ʲl���I��Q�fS8���8�um��(=s�}��!ͤCKHM�UU����u[�@�.c�)e@�&p��l4޲�<rA�D S�е(i�}=ގ��
���;���-/�y�&nɥ`����ä�*cN�I�(~w��PO!�X��Z�EĜ<��c�h0�90�F޳n)mB�ȃ�����$�C,�łqj�E��ޓs�B����:S����s5�)�V
{�<�CdbM��㯷M�Т�E��!�"�=\�6b��")�]��;υ+���a��[U�qq��@}M���w��hmwy��b�&s�&U�yJÅ�d�G�e ��}���>����/&�&�F_�;+\ǴK��r��l�*���쩒4��[��i��a�n!�����_33�ڝ �mݫåw�Ta#\�?�#���2+|����Za�p��&�U�����ì�aKK��)�Jբگ��{���L����c�����2�^� �ӕ	�σ�~u �N�O͹� t�g�Q�RZІ�*]��R�X!�0ɍP7 ��|mQ5(��ߵ{�&D���$��[%��؜���+#�l?��F�>��,�i�i_y,@���[�����v�O7�1���]����ލ�\�Tn̒\��	�M*�fݒ�ښ�">�ވvw|hsoB������#U��+x�U�l�N7��H}�j��XD�L?��$`bu�vf���?I���8��"9S|����k�N�3쑿4j�n��%��.�Ͷ�õ�t��<h8\ϛЄ)��H��!x�+�ަ>u��k|�p��o0*��,��.0�/q�c)4�^�wl���?|�?J��\}�qԱ�mꒇչ�'���
� �2QP�6�3$@x�p� ~F����E�9?�y����:��@\\�"�+��ЁZ�(r+���mJd������OB�c�m>yۢZK��p�Q�[�^�:�n��q1�bТ{�?�-��ʑC�ﱷ ����U&�=�1�V��p��9o�(�5?��qL��ګSSeʻ���?� �p��m�%���/�ث͝���`��	T�[hsĥGx^K��m(��p���b�����(pp��Kt��
�ō�C��ܕ�7\ڱT	eɅ=�l��/a�H�-,ސ����� U�LR���{n�i���+r>�O5�d�w������N^����*F���JL�YF�h X�o��=��K�'�)nU�>)�Y�T@*�e��Ck��h��@vw�Yr���,}�4(B��._�鯵��6�S��?�~�_�OD��K���wc�4W�X���m9w)1A/?qzh2�\@% �|�
i`���l��o�i&�Mx@]����QF���򅆯�k�����*�g�[h�I����u��F?���{��� �W;���Q)�X+Pt?�k5U �m�j���8�C���b�̖`y�3���|r���֠H><� Ӕ8:���q�o����p,�	����^TU�t���y�.Sv˸qT-��!�J#VJ�.���A(L��s���O��5?�_�؀L��6ޣ�%T!ĩ��"�ݕ���0����d����y��[��+��������ײ����K�f��Ҭ�G=���=��[<o���(�6�ɧ���]���L�{�,T% ���+�몖;7/cnb�4Xj�>G>�����UkW~�B�@����Y���չ�m�c���n�JvB��y3�����G�r5d�������9�J�8� uS|8.|�Q�a�Y2���06}��ܣ�>���]O��ۣRt.z-���^js���ɬe�ծm;�a=�3���Y�v��3�7 �,�"#�|������t.��p?��G Bbaa'��OD��h��5�s]^��՘~y���U�c�o��s�����(Ë��F�����H8�3�W�����iJ��#Ю%�`��6���k����N���_c�@�0G[�ũt����(��"�ho��d_nL�|�Ӎ��->�Of��=����}�u�+�}t�v�q�f�dr�B[�!EZ9�jd?��29� :c���=}�I %��E�^���m�%axP�jWم���s"HsK,��+���0�᧵���B3���u�����!T����@l2ѴQ��.�2˪m�B����F9��ԅ+��˳~�4��_{��r��8Mȗ�z�]�*Ɲԃ���I�n���/l���ޅ.�����>w�4>��ֽ�S���2Q��;�*��܀ˬ���qD|���xR�0�Q��2;a�s�#����Ⱥ�w˥�	����vx�x1���ؾ�R��
B��`b���D`8=�$_������ z�1���'�
ك^��RV��ڑ��`;T�D{YN6�%_��QEѪ������"�K���s)�W��o��89�9Y����΅�G |�D��]<:���7l��g8��}�t} [�n����R�#���BO�W�,�}8,꣕$��P�	�K�"��N���&�H~H�	�ԃ��9B,�T�b`��A�������lc�!&�`��؁�ѳRYry l�]������[�Lj����
��{��C��z:�p��7z
gg5 � �չW�4��Ķ{2;!|�)�ҽɦ����5?b(��Z�y���y3ld?��V���3������%F�<ztE�H+�&���>f���b-r�X��s�lq�5ғ=�_ �6r�h����?/�/�X����5��Ȫg��5X���}����nl ���0k���k�p�W{��[=�pw寘y?An�n{�X�K'�6�NY&Csj3�`�N�>��L$][��Ĝ���j�$&ț0�����B� /�]YMF���3(G��zj���,�<}n�㥭aM��`��2`��9���mŐ�: ��!���L�h�a>̈́S���u�=�R]���C��o�$��wE=�- "!��$$e΅�9�m�;��F�Yb���nq8�L"�t��"��Õ�#��!���[/Z�k����2-�������#�#o�` ��2�Q���)�D���	/s`�h�.�9��.��6��^RS���^Xq�PT:}�q��z��^R� K��!�Iz�R�3�e�;�#���C]���S�]���"ߐe)���34���J�J�{�"��.jڈ܆h��y�q��m^ٕ�E"���� ��b���"��n7�X���|��?j�{�~S�Bu󣷧�6)4Tгx� x���VE��I�,��!P��m�l���ĉWrU�X��W,:��ѭ��W�/��ǧ���r�����a�X������"5cK���<-Z��Ph�@����4'%��\7��� 7FQ��#�m������礼�!��|�e/K�6�9�v���:�`����8A}�a���L�$�2�ċ-�B_=�4oy2����Sd���,���o4L�e]��c���81Xƙ�H WW�9�d�_��>�8�q��D�(�?�~����~��Xhv�W`�B�^�34�s4B�����l֏����o����Q=�эD��|��.�ϊ��	�{��]s��0,�R��R�{[X12fkK�o��8�(mƓ�3*�6�d3�՘�U��B�c�-����z|�v����s^�^q�:/���kW���&n�N�l=�`���CI�#��y-�Qdշ͎�q(�C����������t��jB郎`�Py�	�+/�8�_�P��]������BX�yn��s��'S����/U��+��i:�Kr���'���������f��u=�Y3Zҙ��nhE}�#�ٲ��C��+�}`��K�V��U4Gj,�
�tWW%���~�W��F��ST%U�L"��E�����B����w,��S�&Ӈ9�_c��L|��z3P�߹��M1��k�w���2��l�,p<�{���܊(i-��b:Qr���ŭ��.a>���]�4�6� ۩e����u� �?$�BQ ̿^�6�b�qHt%��MZ��t�l�{�$���������Z�R�+!I\b�d&ӧ��Yrg��R�(}���r��t��}�=8���Ͳ����-����|�"��bhN`蛁�bP�ă%f]�r�kk�����S���`*�zL�re59�H�	+Yl��>�!밿?�����o	J��u�r�95J6�#�`��W^hŋ�D���6�`W:)>�4Z&(�t�����CF�����G6��cq~���;P!�ƃ��"�Z��Cj�G��
w�>��h����1~�q�Ϸ�lzl��#�BQ2j�9�*�_u[�)��W�P�[����F��`�	]�\��fnK����ݲ)l����B��|!�>i菣7�V{n�v2T�;@'�g��Y��ump���[L��\�R�Ȓ�M<�|��/�+�2x�V��W����؇u�/�N� �JZNL��;����X���E+U$�������^B����DW�L�}H�����"[�,�'҄R1 ��,�ȖC وL�X��Qe�(e�t/k-����j�m�Ĕ
�p}Ԩ�כ���}d���VbF��������|m���]�G�'J���O38��fUt�J'-�r8����sJK�,�5�-w�Ȟn�OޫL5��̈́O�M��]24[?�0qE$���7�h
���^���~-qd?�z��ƺj5��y�ip��0�x�RU[:Wbb���IzҘ������"����齻4N��g�kU$xx؂�A���to���0t��}t��E&ÊYM��C�Q���jp�jg)�N�!ύ��E4��"���n4q=��3�}=�V�\�0��i]��̃w��i�4�؁+�k�%�  Qjo�ePհ�/4`
9K�I��՛!v��svN[���"*�༛8�P�#�9d����UD���t��m������Z��u/�_(�����ɟ�
�hht#&~,Wc�H�2�`�b�Oj_��"�3�}��	��
�����Ւx�ѡU]Ѿ���٘�А!�]M�<��@�[sϙ�<}��b�R�@|�&�K0f�}.uB��W�u`�5� 6�D �׆ J����Gd=t���>0Ό'�$�〥Y>�3����4����ޥ��t�h���y��E��,�H�L�q9v�nsY�+�'�=���]x�DOsD*Z��@)P��@d#���/��W�9�F��5��F~%ɫ�J4��֪��A�����<�g�ϔ+���4�ۅ�U�1zQVf�Q�luu\qZdzs:0��GdL�Aơg�Ϡ�2v@�5Y���ș�/��sF���� �SP󨉰��'x$Q��T#�*���A$CX��]O�^!/�=k�pZ٣�=PM��B�#(��U����2��I�ɵ�X��"Sq����)��xp}�뱃���^|��p��*��3 7$�!�����Kk}7䚍 �����õ�!�ӀƘZwP=��x]	���k��S؞br���BGىU�0��[{B�U���O��UgA�oC�aLq|}��rۄǔ�;K�S�i���ɩK����6�;�׆�2���������ɋZ���FUub�B��T7W�O�0�2��y���>�m��0���ً`9Ԧ^ �vL:Tm�ރ!HbJ!���&��g�5�ُ䫼�R�77!���h�o����`t�����	2��Q)8џi�֏1s�wP���Ek~�:�T;f��Bf��`���(-r";%�4v��S�^|l�<�0�v3L�DE�.jQ-F��g�7��w�.��	ꋓ��)�&{���Iz��W��hJ��ťe,D�-YQ��Mh�K���t-�����f���������!�,]?�����6�2�&u�w�|�
C���a���R�4^��2��$��u���t����Q�]�w��>�
����ŭ@_Z�wI�_��GkX��>絗���Lg47�_�e�G�;M�\f��|��kLn<�M��(`�����*4��' 	���]F��؞ ���A�!�}��`���P��9�'�ƅ����2J.����>.6��D|��%��ǰyGf�s����˓�����9��'=���Ȇ&!�Z��*j���2?�����U���%zrd�������<����5�gN.Df+|����X+���坣�;�����P����i��)-�x���}@�I`���-����*�iW��~�� w�߶erT�\�����A�&�.�!��I �����~mK)@Q��r�%-��7���t^����&�O#��?�`�~�QU��L�Gg�[4�"���Z{�MO��-���m6ߗa'c�)��kogQ/SI6 [S�%{�$ȇ5��ug[�|#�ˣa{���!%̈�����<��~��w�&<e^/��
�:���I3�ô�)���O)����;�_�5GZ������pvd��A����a�y3@����M1g	rʋ�z�����n�&�>�-��%��T">C��ܓA�%@��;�����M|�Z��nX+�Xi�Z߫{L}X�����$�3�5"p_J���~vྡྷ2�z��O�-؇y ����'��|����zn�u���d�Jb��Y��SJ��zG:۩��}M��T�h_�hm҃�+�O1#�
�9%���jTgh�I�����-���ֆ��b�o��Ne%�@z�1�ZGk�|��%�j}O3���^#��=�.��C��G�s�:���S�!T�i�U�{^ֹ�z�z^Q�2���]z>.,sv|�ў�{�m�xXˆô1�,G~�X�^m��ȶj�oU����nWB�I4_9���~\��+��y������Jfz?��\R�#1^[[ؽG�O�3l��q��g�eG��7�=�n#M
(�?�����ONT� $ގ1���)C�;�����`�=t ��ヴ7L�'�_A����^���:]��,�N��|}k�d(�Gb��Z�ڹ`���aV����+ams>�9ּ��w�#����g�����i�m��b�_���C9I�
-�Aa�[�{Lw=������㓻�h�G��lAo�l�.�$�kF�IF� g�eQ��v�j�B�� ���B5��Vp����
���t��nH�ڽ��uLXސ+#w��ʠ�lȠ�JL`āA������L�%�.�������Cd���g��q��9-�H�e����\���µ#�y�?L��4!)l���J�H(��	�cW�-w)/,�X��,�+���̋O�h��d=�{�ϛG�!,Ȩ��F���u����2��GM9��
��U�ZJ1"a�����'��dPL�����0o�~���Է�a��V5�����@g�K�HE� �L�k�������m)���u	5��5Q�
�P��0��86!�����L����SjY���k��5H�qr��9-�륌��+w׸C 0�J�k������ǝ�z_��k���j��Es} �|��RI��fr'�$�އ�]��ʋ!�����?撿m`Bt�j�Hmo�K�C�%�G�&V셾*�E��V��\Re��a,T��e�9�q�'?򐩲�ϲ����BZ�
�c���������IV<�0P"���}������߽`��}ԙy6N�*%�@����`L���$Z���3<�8U?ٹ���h�	��[dk��WEd�J�ڑ 
[��o%�7~v|�?��0�/��!l�d\|+����	�2�'�0��~���9��HW��[�Ș2����'�����3�'q���;f��q:_9�aD�xǩ���Sp�����D�������Y"�F�� )�t�7^�I"��TI`��u�{#��Gv��lX�^�6͂�}Wn�J:�X��$��KK���$���ř�Y��خ����xR� c��@�����u��M)=�1���nOY�ü���-�~��.M��.[�&�X6�Q/G3��i%vO����Qv֒���G�|!�֗��=�M�� 
�V��/��0M�����	xѼB�h�~Ke؍���	,�h��Lt����p:t��4H��S�^���:�S/�����8���82s�y��`��TG��4ɯ53�.+��ŏ>s����G��(���!hPQ�����4�I͌DY�1�zq>N5H��B�3�k�de�&&(��ճ�kR�]����ɐ5���G{�ը%����M���S�>�kⰀ�.d�"1��5��^ �2�j�M�7/����鲨'����#�v{��Z-v/�_�bX���{F-{Ϊf���q�m`\e��֘�4�.�G�/�f0��Ii�wɏs��'�@����|떱\���o��J���+���m\�"O��F��&�QE��>�
���=x�d�Ti˹X��le�+<�����0��a�M���tY0�o�`����"�A]t�
�v�<1?��ܙ�.�C�������[�#�by���}����@�P���Π��/�� ���ր���k�@ɦvZ�ʴܠyY�S^�p	R���#l8�HM��nZ��֣��@ ��l�\Q7��(���WĞe��4���Xo�?E�����g�L3����̓�<0�H$;���q��Z��9���j!��[a�j���Oc���6=��GI��a俔��{�t�|L�?��~̉~��~��w�n��[�SxGE���=���z���fJ~�EnE���(:#2��뮇%L5ؐ�Č�l�h�]Œ{*�t�,�����*$�lF�J�~s ��r	$�-�N �w�{R�z�E���#�ka��`so4#$�XI1_��&(Fo��?k5���6��O{�-4�n����y��L����Ʉ��`Y�ކw(��r�B7�ع��ͺK��ɯ����/�� w�q��4�A\�����>]�;3�Q�����i����p���� c�]) �>�VBP�`gHL>��O�W�<U����V��X
�G��)eF�'eƧ���x9��A�U�Lz�]��R�q�9/0�[b�B���{��MY�Jp��x۸�j,�P�w��xfn�43{�K�{�M�B03�P���_:�R�ns���D���B�ޮv[��!n�k�l�hD8ۘ�����8 ���c��4b��8^�3��ڬ�ş8�Gyȟ-
������8n����n���������tnO[ùXA�����t'����;M�_2�O��+��1�k�t6�P������up�־�;�$DExig�'��1ԯ5��d��w��K��$�R��>��8f�r5?s��q���X�,$��C��.�ko�L�0�R���b�¦��{`O����X���f7���]��~M�s̅��VSAP����w�Zd$[�.M���1Ao\@ߖ�MB���%�,M˘��n��i谹���Og���J�.ɫ9I����-Cԓ����z��K���1B�
/n]!=��^j <��c�=9��Cnj��Z��ޖ�Sp���y�^i���N���������G��V��C�����H�����d��,�m�v�>��BY݅��і�<O<�J�וmv��2L? �'e��rc�Η��)̓�O��vO���M���n�k��H��)���j!�-]��!�۞�〔x����,��-������s�y(t��K!cH9w]
ɡ��/�[��ou��.�4�b9� �ӟ�$����p�B���W"��>���,D���O�v��jz�Z�*�}~Ԑ��w�b`�TH�K�yKujn��^�@�=��2g���6��`����x�0&F�_YiҪW�}��ӽ�h�=z�m_W���[۱��B��F� ���s-���>��c����?�wpL}���J?��:�����g����F!�H󗾯e�̿C��� ��za5�=��p�4)�i���b��t6Iu%�C��oW
1m[�����~���D4�t�۶%C`��AD�h	3Ӱ�e��T !Im�fi���#?���]k�?��$zt���B���F8�?�/,#7H��ЍP�j2u�Ϲ�td8�yṃ�Sw�G)����J�м��슐B��x�,:d�1�n�ďK%L��s3��>�'�����^(��E�h�e>�`��R��N�9��'K�%��_������3����Y�m����c�)wZ�a��Ƃf��6%�������	ı�{]��D/g�U�ⷾ��T}�r��	��_�\�����'����$��π���jG��t-\M�9t�XR�Al�T������~����3H���6o@ŗ���Ě��Q�_��
&P/2_�j��0����!�W^����Z��Ith�f�(UP��E��^J�U8�P�c�)ɰ��=dpD�g����C���g��&z�l�V���]y�kZ;�y�tc�T��W�����#UU�x��� v��Lč������r	����e��=��39l>��*&y�~s�w���&YJ�S�h�AL�O�a�I�E$��yf�,+�\/��'�I�%W��X򲗦m�<��2��-��-� E�6f���G��a1�xpՀC���b��L��K�/ 
�BxP�Fw�k�����z��Û��ǰk��G���I�o��(�PG�����"z,���~;��,���"���)�.2%u���Ś?n֒�h�����y�n7�[)/$?r���P�m�j�
�c��'%^��T�b"~>y3C,sH�so�.�O��B�~���d���M�:����*i�4�C����(�e_ɦ����5Dr�L;j�.���n��fl`]���z��("IѾ�E��a�хgP��$)�J��y����%��C|aH;/m�%��E��˒���dq�)�={�ng>/������P��u����]��7�9~���;p���s���v��� �o"b�)3_����+$����S��o�'7H�ь	����	�������i��^�-���w I])�� ��t5-xf�lGNc�Q9P��3ln�}%��O�� ��O61�9��<�t~�j\K*
�ǝ�6ٙb�U�J*^{T:��-�h\�C�2d�0/�?��|���O"��E��xȅ�Sq�yo�]�a�Lo.pIՎ�@��7�yx7��Tr(���qջun�fF�����Z��@�ec���Eٓ��1RzCK�^�Z���HB}�a[~�i��|�t�S�}F���FLc��E�0'.�n�u1�j�ȷ�CK�o"6���GV� <��1(�	 U�;���*z�?��s��;"j������%E7q�$Rōu��@>�A�[Z�� /䖣��C&�B�V��/GV�&4�!\T�9dxn�}I:f�Z�����@�#_g|��V�"��5�\�#��N���i�x����ڇ�5���Li 8�mH��6�.�0����67߹\Y���z6�6ޛDR�Y���d���5����WU��5h���#�کŐ�*"��i�o��Gn�B�rWDU]]\����:;x�G�c�S9�}q����|�	��ak���>�ԝa�+�AM���26�o8�VH{�A��`&y��IZ,��ؘ������_?z� ԈE��YEi�F��~A�_�W��
m�*إ=������	[)hA m:\�SLʈշ��O��d�p��s�2�Y���0~�n$^��xJ���Q���T�:d%%w/���t�n���{2S4�s�F�iN+ ���
y_eJ�HS�`���]n�r5�ond�i��=��x	E�c�.�T�%|��~=�wG_sZj��8I��rWa��4!O�kjl-�� S�1�B���R.��tk��E�Leֹ�+���6���lG�F�|Vֶ�n�v����D�)�gt2���1�c�z��YΠ*�B��n���GHΩW��/�t�f�FY[�6F_����೻wMe�ʨ�V��x=��kJ���xڬhl�8���uY�@D$��Bm��k$�U��MFj!wY�~�E�T�}��Ǹ�sS�s�D�3]/r���8&kб�lS��S+��_%�cJ�8k�<�����r�Y� ��������`t�����5C��%��D�g:p �+�a���U�:p�gU_���g`��(v>3�H�N9����_�0�yߏ���:�ΨCp�.׺���D�z���^�z�GO2K�ˣ?��z��u��)���.9�m�O�VH��^Bc����2�8P-Rp/�e�y�ǧl2�2Z�f;���F����E$��]���W������8�"��i0r�6�D�p�)u�������#�SqKk�(G��g�%9���K�P�Q!�X���u�P�H�q�
%CSD��*�Ǯ��t�:X����}.2K�(�'�ΰѣ_�Iv��Y_��_oّ9����胵���XT���^�.�<K��M��� RE͓�u�r����?t�+%]]�2��_>Qk.�����w)9��8ߊb�����t]ES�6/�Pi�4JlS0ܲ���6	6S]�w��4��0P�ph��]8�`��קe�fY�/�C���oh�4���:qB�զ~����,����H����������$>k &�į"o��K���a��æA��֙��0��C���?�7���`IөpM���JY��y�#f2$^� 5�{�.xSQQ��^ы�kVSw6X�9�O3�X��n4���?���C.�T���yD���P8���B�i�5�C�e���Z�6������@�F�b�<���ۏ�U�ݥ݉;���_��)Qc��d!=���S������M��j]tL���ƣ��C��ʥ�X�K��������]#{�������C��DR�=����	M����}=��g{NFyK�R�-��w::��;����sFYJ�����H�� �\�>��o��f�DʅK��&��u��K�2%Ca��n=�K�ξ/q�p�`zQ�
�r�K݌'�����rH�SB�2g-;N� �2s<%�=�l�Ӯk�ee ���^ �I�jj"����tYf�4�.�Ws�,d֔�0]�E(�c ���Q+p�!8 ���v
d(�xR�6��)osW�(�P��&�H�A�}c��,����o�7٫�V������\K�j �tn׃|:>�<�݃0HJй_�Uݪw^�"�b����4m%J��6d�}���R�3��?��T�N
E�j�8?��#)�838\El sV ��2!���L��޸�*&�Wnջ
!�;�W��íGAY�)�������AIf�����h���L��2���Y��N2M;��iK}=��@�e���2�-��Y.����~I�m�h��`_���Dt�2�􀍩�Ԋ%m�:
�ԛ|�*�1�("{r���WCX��Z��뛆�'���2�k���N���(���ƶh�V�	��NҳQӢF�$�p�YL�Óÿ��"T�K�N2H�L'�n��MGV�t�B����p�v���v�V@�`�(�ۺV����Y����y��:�� ��֐ZE`%3S� �v7��G'ӑ�]O�A,@#�c�����n���m>����8��+����ώ�/�q�^*����I�,+��j^����ﶾR�>��ƕ �po�"�:b�z�*�h�ٵV���(*���.�MM�&7�ƻ�<������1wVr�b��Ak�tr����P�ʉ�^���QYk:��y)Y�m�1?_�9G�7�e�2���=h<-��QE���b}�}(㥼	l,R�]� �v�&H�1�t��:)�[�߹�v۸�
��T�VIs�7��l/l5�b�]fF
��\Z �Y�&�B��d�PO�9=�E�+��<�ă.��V�ɯ+
�G*����A��Ư��!�m�ce����b}����g/|f�0�a�܎FLa�G��=+�#j�	s��/xi<�)��/0Rb:����(���ZGׅ���N�ē?| f[�`5,=i����_��o��wt[�[��P�q}"���=Ŀ�Oh����H"WcH64���Os����`"����)21՛������=R��
O���(J���DU������� ���� �ʇ;}�R��8�^[�}���Y���<�jR1T�nΛc sP?�;�=�qn
�n�'{ ��b�^ERk���|Sm<	�fZ��z�/3�N�X7e��rqV�T��j�y��hN�;���p�b�ʟm���������-΃�x�yK�������/�3�+�d:�e�1胄�$说B�gd��5`���b�e�~�.����S	r(Kl]�^�a-Z�1�V��逵��z�j�vc���(��W�p����"F�?#4��D�d��	|V�_�(���ͿQʐ�J�Xy9��w���LS	f���"�IS�҈{m��9W�W����qoV=l=��/B<F�"ֈ͹�X~7k�.&^��]r��l�9�
H���۬�={z�w�fa��n���	Tp�ؒ|ע�u��A��+���!y綧ɗzI_���A�sٱcB D��-=�n^�E!2����f�lmuu݁\��lzN�I-H-���_oM���Ts�Ҷ/�K�%��U,�,��Re�4���"���el�^���'�Ē����
��O%Ңt��[3���J��|r;rM�5��Rȇ9�� �!���]�lQ���::�R�!J6�>o6.��o�Ws��;�.ǜ~��.���:��Mtk�m���ۏLp���?�-�j��f��ql74+�aH�"X�Op�𖹶�{ɡ{߿����z�8.m�������܂ob7���`��u�6�!p�3�SH���L��BsN�U⠆)��HB��C���<l-�h�molxN�vkz����h�10#