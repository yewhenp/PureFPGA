��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� }~�XVӕ�4�3Mn[��n�o]9����ڮgS��w�rB�^�*�'���$aX�x> ���Lo�S� �,�)�]ѧ-�L�sh�4	�^j6�t�ͅ�>@�I��:e��١�E��]���+�)� qц}ad`�h$>x�+��Ri,�}�U�sÙ)n�!���yiq>��ځOD�e���~��0hKf���U����;n�U�CJ�����Nx�Ⓡ+׻M����3�(;U0��:+�(ީT�#��g�4!(��S�be$�p����,�w|�E8㉅������u��p���)�N��	�]t�:��f��+!1�{P��0���ɨ�؇�Q=�Eʒ��V�*Y��~��vs0TJ�Iҽ}�s���u8:ɖK����rl8��L�!w�E%q*�f�#��5�Kq��ۢ��!�$3eCo!�d?�i���~�*�m'㳣r&��^ؤyC&���X�,H����z�I;�i��4[��D�ދ�5�@���rdӥye����Ti�m�WJ��"��)3
C���/��*��1Dy����X��*�j=-����%���v���YΖz�lTA�2��Q�h�Usn���@����n�}n�~`�5����x��b�^�5Ϊ�D �DKS�}��N��$j����Ɨ���jI����!���K	*��ڣ
Ά�?��mh� �=͓%�)aj�ʛm���
�NB�x�=7G4�MZ����u�2%F��ΡĘ���=S6�JDW��(�����:7�c<A������5��*S���VV%L��Hs���0!8�,֪#��~��bU���"nQ����V�-���8������L�_l�<3D0�0��~���2u�p��ط
�;hАm�f֗)Ʊa�P�QT���^����/�q�;?X�QZ	cM�X� �(O��V{Vw�l�j�P�i+#�M#D'�v�Q�n:�"t�(��<��x2�`�k��'h8FL��-$E�F8�В�I���i���X�@S���5�2m�!4�?59���Fq?[ �a�I/Ɉ�	6��������%���i�f�c>��������qi��}�q���Ӟ�9��]/2�����+��'+c�qv3!�],Z�����ܓ�1�D��V�0� b�8:g}y�E0���[*�6�d�P����5�-��U{��u��-Q�q(R��5��7�-\8��`rkXK�3zO�G�<O�0�ļ�Oz�dB ��Ӻ�q��@lU�|�bY d�%��:�1�}��b� ���<*�אU/ x����`j� ��;n�"E� �8z�bxd@�A��V09R�!� (�Hw��e��v_?hy�� ֯v�"����~P�t(ӟDA5:BP�Ջвb�\5[&$�Ņb�f�l��z_0�Sϧ1�ªܕ��z=��;FhI/�Pv��	$<�|�%�����4f�!?��x�C�A��e����4��� !���]-��KM������1�����
��Jů�}� ����b7sl/,�Sӝ�7�f�^[��6%3�v0�Cp$�S{�԰�_rb��'�w�@'��E�ځ͍-��yg�Qg�J�aq@����F����Τ�t*<���}=`��ds6�U�{�B��- �p�.<J=uI�,=~v���}��L��@qt+���W5p�s���3���8��?y]�:�	�3��?�(2s//�*��v���2���Ɖ�{��P �:�7O��_�E�v���1^eC6"�Iv����}�'�e^��7���o�O��������H�n`�2�T<Z�����E:��K�)'_��4 �9���(c������2��z*��x��%JC���M�{rʷ_`RM9��
��J� �?���/&aH(u�Z�:��lzd�9hG;�s�+�o����yT��c�H�/���)dJ|��U��=\�4 <i0(Z��| m˃&V�;��kW�g�	���s�gizp�I�k|샢;��LY=ZVE>~w;0�T�)�}��n�%���,Y?L���V����w��f�m�w�k/�K���E�Jn︄��� l3�����+a�B�� kQ;����[�� ���{�Q{���"�W�Ҫ��J����	~Yk����"'-Dy�Uc�_4��ˬ��(�CF}�۰��=pݚ���Wk[J�G�D�D��^�
��n@�NVƽ��i��bv��[�Et-2M���\;H�q��H����	����wD�(u���H�@p�]��!o����e'c�=ޗX�0F �72#�1L�W���B�b�r.���i�`n�]�H����H�h�Dy�IFԜdGؚވ*1䦍VR�.;#�"^)&]ӭ��K:˼�z��z)�ެq��	�EtA?�Gh��`���LS�����x?pww��{
ek�e�q��1��I�"�l�q�N�n��q��Q*k{/��^�����B׃\��9�:fpT��;ĕ����wƽ���Mv�j*FG���
���hef�6�>�#�$Лxo���}���ekV��t.X��J7j|�jݺ�d�9Z����1`]Z��q��P�&�8h)�Iq&߽�?�U �x�(s��p;Z��\T�[��Ǖ�)k�u�9��])�݂�3#�Lm�S����5f� �5Cr�8�<{�Ў/��M�m�s�|I���.�v�1 '#�W��E�� �ߎ���RG��uڐS��~�{�z�=�0Fr(ߌl��T��X�
xB̰Ў�	�S ʩ/QW�K�zv�&< q�aY��H�7<g��"A�=Z��I�s! ��l��q�e�(p��{�ş/3�i��d\˸��=u���zM���Y8vV�g�[�F0���n!F�������w��i&��m��n%:jYLc&TG�J".��`Ws|g�����c��)�QgnIPS��B�E������|<��A�dڛ��K�0x��4�Ғ��<��h�7&9�7O�?��u����b?nQ�;-S�W�aa�4گT1\��q	��?�����W;��4&� 8��S9o�A��I"':���k��?+M���%���7Y�:�d�$�T}π�ҹ#�Rd��鿻�����$�p�0�R뮖��$b+�Ȁ>y�2/�B=W�|V��:[C����]� ��;
��&�U\���Y��ߴ!�7�|�Ղܤ��Z�yW2�։�!��(��M���:�B� <Q�n��A�j5܉�w�t�$���-���rZ��5�%�%o7�#�;P��2��\��T~-���S�^���Pg�*�S��T�L��̿��;��4c���Y������<B*�ì�[ �y�)��R��UF6=�y$ں��/d�;�L�`WNKn��������u���)���J��1\����!	���~��>��a�E\=m>H��L���iA�A��k�m\\�S��=	�T~�����,Y6]�s�������)�\H,�(`�G����{P�%�P2��.��d�[����jb4��n
S�ak�~�4eSWԓ?��r�G�0��{d�n����J0m��_۞ZF9����V����6gOu�s���4k�,�M8'ҍ���t9�!�@ ���UV�S9O�o�J�#��B���j����zl� X*f�IBS\���^'~d�r����͘T^R�x8�F.�P;�z`������+Q	[}ܛ�l;��n�8�Ck��z�б�Q��N`o%QG�O��{�i�P��z걃�D�y��ڴWf�h�d��"���>;�P
 �-y�`M䇲�`���PxVt���ڳ��ć�ӰWl���.�yF�#B@j���k�J2@��Q���5����?W_G��]�{ެ{��@ ]�2���"��t�1k��A泽{[�}%T�˂�R�vVQ*-;g�+�=��Hv&Y^og&�>���p����=EТ:E����gM�ٱ��t�=�D
o�-�aF-���㩀ܢd�3[�F�R�f�C�%o������n�J�S�׶0q�"�g��>��J_�HH����8���5*	GGT��kS2 O�V]Pj7�9ϒ+�y��f��r�t�"��IBq�ޜ>E�pI�k��m&��N�^����q ���
���#���Wk
�=r�	mb����ȝ�e�ͨZj�2^cǟ ��u�j����7lF:���*\�u�)��"VP���1��6.�.]?7̉C�z������y(G�®���fz���fds{�v[�P��G�#�!`���jCX�������[��M��z�c�9o�9k6�o��+��r� �5����i}ԜE��	������'�jQ��գ��.U�u=H�Co�\+��BC�w:�*�! ��E��;VJ��� ��H�R�u�7e��Ǚ�oG�xҘ�n]_�MÙ
8$-i3	 �@��s���U�IK�cjX|-K����x>���^�Ox�M&��+���`RP����y�����l���-d\!��+��՞���he�tr��6��Hd���3��xSI���+Fe+� ���b���^�ڤ�Q� ���Z���u��N���������͡��l4M��;��
�3�91��M�}�w��?���]թ-�p5�7�mI�Lz��h2f ���� :݁���M���;���-
m&稍�u�f���:*o�N��׉���9��c�]�{-z+�Hz�/ol�x�hiH���4;m�_[V�`� �����#��&����W�P�|�q�0-��S�y���\ޔy�v����靖�4��ͬ�u��N=�#c���[��,&P�kB��έ�0���{L�d>י�p�T�⻙���:��wN��h3��rRN�M��p�GB@ҏCi�[�}n{���-t�<D(<�T�C7ˉ��R���23�(S1Y�,Yi����m�9�l��F����V�@<Wv�`.�8�#5U�T�(�Dw
�m��6�r����H~�q�Ӹ�WX�D��Q%����8(Dʂrw�
,C�Z�#">��oK��5B���F�J�퀰/�����3�3����&��1f�|`��]1v�s��oxSmZ���f�4� F�\0���J���Oߕ�:����e�zg]V�Ģ�6�k�Y�=쭩
��N�
0����$}Â(�="�z\`�t��|k��l���H��|U�ų���F>�9{96O��$Ew�����w���Ǟd��5͆������\b]�e�F0\���v�;���2�D�� ~�Fl/�hQ�ߒ"�},a�,9:ӻ#@�����i��{�(��];� ��O`ڛ���Ǉ���ZR�Z��U������!��O�pwv/�0H6)�R�M�Y�i诇�P�&��P��.h�]����"����'Bu�% m6wt�����%��-{<�-����+��l�[��XH����� �|<�DlqE�v+؅���)-�H@����D{��`iƊ�NR\ƓR����n�Vа�&6�|zQ�q����'P�������p�2�_f���{b�	�k
�������UY�dQŐP����9�r�L��������\��,���f�j��<��БK��H��~\d�h�SR#���}������$�����˻/a���e:$��~��>#��w�sG���\��>c':�(mA��X��2�-n�kLo���Z90�if,2*���E��ӝD�,�-�~��i%G��:T��ل�Ԩ��,9Rwa�.�ݣ�/�ѵ�%
�u�׼o�9��E[���{C"2�O�贖f�tg��-� ;�c&z+6�惥�6�̱@��B�0���x/�z��{_(�'=�W/�Q���]���A�b�-\��� e��/����	K���3�3�&���۞��=3L,��0 _?"�H�)-��4���/,M��H:��e��#�4��4E���9�A��/9ǿ�>I.?�m�q��VX���Ub[k����lI����A��jҨ���UyK�Q�HC~*�}�!���b��)�=.���ۧS++6rV��:4�E��b�;���w�V��KK��ҥ�U�E�O��(i���~^�g�d����}?Z8�1,�f��,͔����<Y����TF�D����A��x		A��pT�玛��)(��Si��ކ�)t<�[	,��ԉ�e����?Q�����O�^��l괒=�9j�{��m4�4g]�ʻ���+M���M��{o�|����4	=3���C�q��A33�Oo�؀�W�bLq�õ`����־��E����e6T`�������>��+gBfL�d�x`Y��� ��s0~�1�_4��
A�E5��[3�}�I��>'����b��t��z|_��<3٫��;�,'�恭������;�j�g�E_4f]�z��;��U�ͨ�g*!�9*3yK��0wdX�XP߰��1��F�N�.Sˣe�-�%�����|��$�x�\�l�4����[����#1���2i�sbs��0%�M��r�lC�SH���H<�U��9&_�GP4�]?�����0��8-��w�i>��1-�d�z���g䊦�ۏ�Z�1��F�%'qv�Nw�F����i#�@\�ԧ����N4��v��Z����ށd�?�D*�`Ԧj�K�����Vk���l��fp�WN+~#�嚗fH�;��ۙ��9�#�Vό��,�wu��Yc�W��ֿ�"���2�q0ٖMR4"q���Gmd��g�%��l���]�:���%$+}���)����f}��(�71,G>�`��||HF���$�=�[p�6F�Ӫa��I1C��QE*�����U�Fiu %�����%,���B@�EC��D�)�b�~�Rw�o���6#%��{(<%t.�ڪ�:��F�����C���Yr�/�[�'E�J�ǳ+���R����e�������_ck���?���V�׭�r ����a�o�W)��9!�*kKڀ|��2��s��6 W���z.���s�ϖ�^���d1�M�2~S�v�n�F�}a�鴑9*՟�2ȫ�D�v{���)��?h�߀���oeϽ7��̪�5�U.>�"Z�I�Mp*+�m���J���-7�@�q�����g�E�����FAQd��Aw�{�ӈ����&y���������3�@��y#��b�T��Ǎ ���n\�h�XJ��1�����ی��?���k��������6��,��Aa���8�D�Yk��ˊR��"��2,4�����kٿ�����=k�i�T=!C��H���ni_n�a���p@O�ڦ�m��m�L��g0���af�L���xܓ)�-r�s^crdv�" fw`Oi�{���OP�������X]_i(B����e��7�}W������9YqE�]W7	������y$}���aF��Q7e�;���𓤝��ˎ��c�J�ۢ ����1ʏ�C�B�g�N�`m�R���$w$f΢Be|�Jb��,�R�\���7����d�P�Sz���0Wޚ�o���d���C8(�i����ũw��i�.+mK�߸E�ɼcE�愋�x/�4�>F���{qh�s�&*���1�7{�f����u����H��qF3a��מ����� ��߱�)��cŒ�̝�j���{DYl�E��:gf{�Z���B�M<D"�R��/����m��mgle7 IU��S�^7�!�n�Rĺ�
���)��-~�`���f�+��Q���H�)�d}^�p�1Gj� 4y�XB�o���ș�ϧ�q�9Xla�nc���0�m����dCB����"�s�l6b �9+�H�	C}@��M/���G欿W�D}�ޙ��C�YR�	f���#ahl��R�ɴ�2�mז�|�1�1��8��-�b\:"�F��xa��͞U���,ς��&`!��ˤ�CA��Mh����P��̛�X~G��̳��X?�H�ijt���{)�����Zc��G���I�yÞ�R�N��`k�M}�^��l�F�Ԏ�;fF9͐$z)��;�Bzc���w����{c�"Խ���됗�~�g�kKQ���P5t�<��S0g����؊����w�d�����&��J�LT���}�)Z�1���4��l���0�)T�<C����Z$ r�)|���Nrix��!�3�<ތ:��'9k�U]~��WD�O�g�A��S�Ø�f����X���Uɿ�� P�Υ�F|���Ъ!��*�Q�6�ȱRإi?��H�{S[-���H-�C�c^� 	O�"MH�<Zog�[�$ ���z�Q�?��Ȇwu] ��ܡJ��`�*�}���i��U߃kȧ�E�|<�����*
ӈ��?�GJwc:����X�����b��G\�h��x1:�`@��ը<�o��NYA�!��}���WrT�����JO|iܛ�Yq��E���q�l"���#0p�^�G�ڨ�<�Z~�k=6	���V�@"�@,�Y�JD԰X1Bv��r{@������1�.|�����0v��J�i�����t�%k"p�V����@�O>8�mS/�7�Δͣ�iI����}4#�/T/z=��j�