��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ`T�}�w7�ɴ��劂���n�T-���*Q@$R�Q���j��g����8�{�6<��O}]wWKȎE�Y����ю���^Y�#u��m�1;�8��Ph���Ƌn}O`���������,��El��C�W��
:���?�S�3M�Ȋ��*P�m�]��k��U ?l�@P3��~�#�;��Y\Mx��,�?�]���9x$T1nЍi�)���<�v��'�=x�P�s�H�6[�{��.a���3�K-F�a65�]u]t߄�i��������v�|q>�+��3��_ F\#���Nr�N�<�Y����m5r߂�3�\/c?�o��+/�B�{�T�ɥ�a,�1�:ov�8 ʵ���}�ola���u|2s��j�%������6��J���F�a�k�x��hQ� �v��ɫ�G	+Ü���������{H�2˼-j�p�I.#��BoAjO�g�/�Q�w�a�<�{�ܭ��'���G�/<|�;���a�9j-� 7`w��y���z�._��=4^��{,�>L�a~@�Y�������	�W�+2�Ն~�1|����	�8-e�E@�b�+J8V昘g7�m^�	��?����+F���\�$uF,�Ps�.(�ӌ��IB��ڱ�=H:L��M ^{�ٯ���SL#\)�j�ܒ�C̊	h���V�+
��
艧�5�@���2"{$J�y#U1��iՈ�08��0��L���r����3��a87򶜯,ڠK���:�����*l7�`o 3Lެ�y�Y~T"�:ʎ[��o<L&w�Ƨ;���F�x��F^;�)*�Je��*n��<�H��ʫ��BWfDa`^�x�4�Y7ly�~���7�	1�ό���O]��I�����;��(DX�0��צ/kC��U >u�1QF�)geo���GÞO#Y��~�Iͅ��>��xpq�ӍY��!4��uC*�ߪԫ+O��62jQday΁ ��@�,����f��!B0qJ�a�.	ް.�B3���}b_3����D|4��]�C���𣈠bx�T87ʕ2����9Qva�H���T�G��DX{S6K�N�l�~9�a���� ����ɉ(I���ߣ�D�d3��6��䭵Җ�kU)��|�}f��ȳ"k�`��3��{Q���,_[bI�c�p��-ӂs?C�u_@x��ف⿺�#<���|������lH��i��2����"�H�E���-�H�̓���ƪ�-8Ϻ?�t�=mݑ�U笜�o�`,��e�V�������y�1Ԣ�'&('����q�_��V{��{��.Z(�f-��쀍�j+��0R�f�q=4�(X'+5�'�G�ǘH�s�{:�Ǿ:�m�GD�e����Oc�X�o�j�FVܔ�sa#�FV��4�Ī���nV������MZ��7ɋ6b��x����/Ve����Qa�er�?��0���ۡ�K����o��M|�E����ZD #�+%�[���iT]�h��AZ���Z|f�r���KW��nR�s�73���Q�:"0 �٪4r[H_�/��շV)�&b|�U��b��ĳ��f�T��"cm��z.���U޴?����Fs���k�[ğm�����<�J��f,�ߣ�!Tb��|��G�c|���/L1���"��ϲ�<$c�KB�`��0Qױ��K�x���ך��P��jx�����F�U^��b��	�l2!;�����g&>틾p�n�h�����9M���˨�_]H@i!<��L#�~p "��Oˇ�6*����$~:�$�M��ZYV�FO�)V2;>�^Z3��WPq�b0	���_�����uj�~�z�y{����(�M�xz��>aq�=�����vl��"-K`��O����*t{ѽ�]찒8��ѓ�v��(��,/Z��k��8MN.@�<e�ڿc��9���Я�fk��[%�
�d�]��GR {��O���+ø��Pm"�W�m�r�L]Tm� S<��$"t�����lQL`«L���j��^�X2���4�!y�{���Gĝ9�*Ӧ��;��&�@}5��t���n���*d���H~b�nG��U�:W�r5>P������B�6��䉅#��`ey�ԏ��Ǣ���^r���<'܍=�������gh�k_���r����Z�N��	�0������T]�Ȕ!�@Wx��#,���4����L"�Y�y��p�$Q��-*%��r��^Jgt�^�g!��E\�W���`�0LVͷI
���7���G�� �pv�G�J��}�b&3B��x�k{�����*�<
w߉\)�^���U[ca��|�Zp��uN|~�]u�q�O�
M��$���~���_wv�qҭb��z_\�6&P�w ��<��u��ߢ�����6���q�-=)d�c�c�	��.2�	%O�CUMQ�Ӣ¨��K��o�Y�y$5yj]	uM&���U�I�k�6U�m���{6�ɥ�.G��𶍡�tk^��i|�������HF+1(&!��<�!q>�`�1a3�\]3:G��Z&ۯ]�/W�6�x���3� �#!���S��2^_��f�Ʋ�k�_�>�(؀.6�;�JT����|W��ٰ��Up"�n|E��Tx�<�~��]?4!�(�Yr��{LЅd��3������hRF<ɤh�_�d�]ُ,W�Hηw�c ʀ}�\�#6-n	����!�-�W�'�CV�������+�99�\iq�|�֫)(�F*%/����ч_��n2�z�Q{"*��t����J���V�M������)�z.��.�5�BX���u���):����4��/'�1)�㌥3��210i����-��xߩ�,�xl<�+��?�z��g�p��W�(��c�S(�)`�G���H��[�G�����&h}`.���9�^٦��c�'{���$�W�����S�1z�?C ���';۞���ij+�:a�K㮚Z����X��U�=P�xe>��S�:�Z�&��qx�&�0���lp
�Z%�� �|��$36��=E�EM��@:��G����5f���0��B¯����Eޔ��If_�o��w�c�O7��-���ۊ�Rp�u�C����*�'�Ǵo<���9*Aq
�cToqJ�.�����ZA��C�8r���u9VH�^"O�a�t�]�<����m���|��'f��eð���>�ǭ������hbh�@��m~h�rbP�bKݧ~UNp���?��׭�Ժ�3���8�o*k�$Ҩ5�E�z�G�M_Рr2ju��;��u�ZҰN*ll�"�)�=��T��-70ʶF�jy�d6v�@�Yw1��#C� r�~
g�D�ܕr�tP��?�4]��>=h?�X��Z��^݅��5��<�:�Q���ə���,G({(z��V���=��p ��>�&��[y��edh�y3!�/w�	�V�_��;T�8�ŭ�m]p8�"�g;�3�sF�:@�i�06R�XB�/�Y��m&�i��E�`�ƱS�����FD��'ڲ��]6�(�<��FOfۍVG���x���8�p��g�??0q��9W�j��!�N�F.�)Y����8Z�Y|���\<��;���*�r[��,B %�ּ)Ӌy����������E�F����4n+ݿ��p,���QH�|���ҹW���DxM���S���6�}\���!�p�ƙ�/WZ�Ӈ���ڜ�5��� �2�V�qC2� 8!w��q�"`��?����!����]�����x��ÆD
������AX 3�K*6oϣ����g��>��FxeA��R�k@�E�Ĭ�b��&��Eӳ�&��u�|�=G��!֦sB譩s�>�B�z<�l����q�h����%]�h �崱]�p���??�'����4JX0	�4��z�O-�?ԫ����TJ`��D�����O���c��k�9�R�Q{i��Ԍ�W��tr�!��|�Ӷ�����*�q�OC�!���i����D��$�eo�(�ݜV9�G�\����̌n$��	Gʟza�Sj�u|I=��������� ��č�0��/�_1T�WN�::�_�|s%���j"�k��)<�ކ��1�����+�1�$4B�����'[_�T��<�ŢO�;8�s�yl��i������Ǫ���˹�Sm�;��?����k��'��P�ɐI��g�?�Ojvkvf���^a!)� �ll���@:�V^@J�߻�z�Y&�����u)K� �;��g��a����?L���.G^0K\�K*K
���d�p���]N���]�e�+6�1��lV���s�O��w߯K�y�
��@�fG�{%�	����G5���dn�2�)y����RD���Cj��\��K�=X@U�"C`0�	/{��CV��iK�5��T���1!�����i,���.v57���0I;�D��6Zk��f��A�^Y�>����wE|�>��G3ןh`�h��1�����)c
]ِ�:�~���k�׮����=3���T���X��\��oݿl'���1-/��yJp��$�O�,ȿ�EH(1��܇�'�!)`���ų�_j���NS>���͒��il{D9r�2XFx͟+��y|}�NnP�m+V�+%�݉tb��8���� a+g�n�0����X�O�� �kg�����v��<}-ղTg�
�#�� c�\S9H�Ӊ�^�ߘ�lbl��������V��"�!�8@8:�˛XpOr�>#7�\�]� ����ǘ�ѫ���r����G' �gG�a���o@,-��
:���G%0�M=�C~�	�e��b����qd�&���+!|=�퍦:�~_7���C��^͓�^O��ʟF���8��v~�
ܯ�+���솯iZ�(�߸*n8��_ֽ�T�S�|3\��F5sMYD��r��M�b��̩����\����Am��W���O!�o��S}
�=Pe9��X)^/�E���w�����;GK�ac^0�,Y�:����&�W���p���=�aL�#{qn���y ��rb-����(:� ��o�:A�z`��h��i���(��&$C+P�tKJS�j���C
��-�{�&�)9��Ni��~�Ȑ�BI����*�Z����aEM��q�d/��ĺ�D�Q�t�nZ0�lt��aյ7E`B���q�%şu8y�ۂ��0K���.�3���Q���
b;HC�?D��5Y]%���� oO�������-3s�5k��YE�ǅ:�Hh�IY��~(�yY(��}h@�"zDѪ�xg�C�Y�,׼4����A�,@���:���o'�vNϖP�&U�������L��W�������ޔ��η?:5�AЇ��˃���@�=i:_w����AW�^A�@1c�&�/*��p,�����*N��;��θȧ�bP�W72�2_%�j�{I�˂���g	����m̹����5&䙓u���©=�(�f-�#�;[Ԧ�`a�!��ʟkj�Z��W5�P�W0EX�#��J[ ���-y�3]�L�f���"�	��7�E�	+L�e*Q�{��:��u�1����χ�Ш��^H`M"�5�p�T�� /-���W���=5�Z�=�A�;|3j����9��ilU׮ͨ�)3��&�C��S����� �}g�%ƆV��W����ff�6#ý�i�O�;�D�N���`���H�d���zأ�ʖ<uB6�R�Թ����>���8���+*@q�A���ނ��0r�;@�w0���%?�f�3���Mw$��]����T#!�g)��pO�$�5W����d���qz�2�7�~������F�Ⱥ�H�1�Osw�����3L��c���ڮ��o���H��ɯC��Rl����/Y���d�xq�dBy?Z)���ps�6�}��=O_�2��m��0�ӄ�vAx���I|�tk����$��ErZ�f~_~�V7:��K�/!�rMbss��ޮgU���¬����~����F�s9��2	��F����0ݿ�:m��\c��M�'�]�@n�D�qCTc�,C��2�9�6�\v�R�����*,�dlV�̀*h���L➛j�8�v��b���oc��A{حXg�+o�U�U>���y����r�E�g��hdJH�12����)8��5ߕ���Ţ �R��;K���&������t��u���=w8�bh�H}�P~L{.�7$��c���?Z�nE��ލL��)]�i�B4b#7:�eܩ���G�4�܅��hS��{���K����|����8C��v�=B�?��h^{�����I��F��jK��#U8���\���e�t�	&��Sح�!&E��rz�I'C0c�����|~検���/�!a��	�>�'U�M�%�w��Ǎ8�������o!om�4�	�,��'s@5��j~9�T$��������]D1�lU"� �`VrDp�$4��D�.�r�ެ3���ڷ�LC)1�W�ns��+b!����m�*2.�È�u�"Su�v��Rl~,�5�mi˵�!3^��N��0��`�1���@��ؙG���mw
TH]4�4H���lx�ƘVz-F��k`qB��3.��h�EE�ـ ��R��+ԫ8���������	�

$�EVfߦ�h߾%]��`�V�ڎ�&�y�@��
ր�3d�N{�en�Fo�r�2�4'>�Q�+�)�ǞA��cR1i� �L���Zc΢]�W+��N�|�c )�6���W�q#�� ]{�J����ոi|��G�j�v�|G�MY�Ej>P�?_�x�)��"xDb"zY��Zu&����x�&ȼ�5#=�YL�P��A�0|�T�}���&����:�5"@�-L��GKK�ɠsD�:��u�<�5�J�*������6���|�Z����6.�����Jf��DVܳ	v}��Ł�{|�bK0!Ӽ���_�r�I�T$ڈ�R��W�k��r/��⤯;�W����d�D�n�&4�3-+L����D-������A���FFäA�m�o�8�;��6��A�XA�Cd�뢢�Sh�Em�,���
�2h���J��p�~J�2�|�\B��\.́4-�I�~���gu� ��$����yP���x΂�D�9������l6���V�����TM���{r�E�k�trf�_��l[]��+ޫ�`�H�0��E��G���~�ʦ��Yh����7�;�z��#�}�8�&��f�K��G���x�:ڴ�o���/t80���[3�Z�`	a�`����|/�K���HY��������}�]W�\��n��`��?<�b���[���7�G%!-E�i].�$AU��N����v7��
{��g���q{P����`�m�/���*��=L�⤁j���*�hu����#��y� RT�*��6��RM�`�+(�Pj��������5� :T��i�Oz`bß�٢��f��j�������=.Aؕ�lK`>�T�1#a8ɨ����tY��O��.䘒B3B]~�[6�&�8u՘���h5�x%��G"��2� �ÿ��_�[�3��P$���R����Z_��|�N�9�9=	g؃N�'�^yĘwWg*��̮����Kj���qK!�\L��;�|�~�g�_��.Y26��F�c7rj}���Gzw�R���#�3V�o�t���K���pYz�zY�Τ��v����t��_�ē�ɰ�ר�*4̎+5?����ʽ�x�r�k�@>�R�5�-$F�_����k��2۳R��}�cȇrp�����S�ͺ�r'>:c]B\�=�F�z��e=�6���V%��Y�X����<n��݅����!���G��R�E�l�!���C(��������E�k�����l�w`ܑ~�.k9��u`Q�R^��D�
�r��VM��f�-G֛��*�� �#���;k��r�����4k����G@�b,��=m�莚@�V����57*��wս�к�A7�]4��~���|F��0�2�M�r��
	H���k�U`��� �^�=�!�-�0�x	���wR��V�t�p*��9+1h�6ρc��;� I>�;0D�*w2,iTu�9xO`p)���E%{Ӊ���.�Bgm��1���J+%���O5Zf��ա4�R��4���牊�8\��K�������GQ��Wh��<�Z�6��IHZ� ��Y��|��D|�9(&o��R��qv��w�ƣ۬� � ��2�Y�j�r������
*���z`��7e�3j@�����W���!�pS5ޟE�ڒ�4xB��AZbmE��7}7��m9J`�����(>��^�&z����P_��'�=@~�tme�_��Q�U���3�q'Jhd^��X��*R�,և�31eq\����]�ufׂ��`5�T�m�n�����僟�WT{�F�_qv��]�����RS<��n�3d3٥k����˩���7K3 wx����y���r����B��K�]ld'�e�R���S�����Qgv���߽W�T ����p����:n@lp�%����}�1=͘��8`d�?`���=i�[�i�R��B7HVE�1�S~�;�Ķ���u��xGC㶑yՐ)�0���X)�/��}a��2Rl@ �W��c����ʹ���������]}w��~�������1z� %�D��Wͷnm�5,� ���u�N^��1����O#�����Vo�
>�N��N�Ae������L�,�F�V�k
(#|w � �Vˠ%�|�.Bw2A�&#�v���,c�0�@ゥ��V�C� [��	~ƭe��lc���/csr$�7ۯ�dUE�����ϋ���ܕ������.w´PJ'�49�0WQ�S���2�s���f�����5O���D,]��Ƨv�I�_[��#RL��LPn���� ���0k�*ھ9!H�]
0~����"�(��+f�޽������^T0���9+��N���Z�eE��Ȃ����!S 	AGv��^�HE,��>i` �m�K	�L͠XC�,p�u�u���|`|1Y6�Z��].ڃ_5%3�0�'qY�<�;2�Wll�(��Y��R��ݫ;�$I�<�^�zH�l����}�8�����2��06SOC�a������H9�vk���2��,4�i�h� �zHç����?��r�V\�C0�xZ䑮��0cr%�݇��^������D���:���)���-+䠽�Ln�;�^t#	�F��%[ƾ�]��m���s�7<����f�v�̹U)~1�J>7�ԻX�R��� o}W2O4��#���T�����Qb [ ;bvǄ2���*}<+���Syߤ�B�S�
lm�n���1��M P@���ٮ�DEgx8݅=���!}�9�ԹO�z���;���h��GX�w��oC�i�#��	�a�A��X�yʹ�Էw��7�������+��M����ˁ���UжJc�7df��s�/(hQ$g[ʏKY��p@P�_�קX�b���d_�?�Ʈ��|�XDp�R	��RS�L{B�3�N�N3�J��B��eb���c�����������~��q�Q"�P$�lI�m-z܃I�D�Cs�꫽r.�&�)�IR'���|��%�߈0a��*g%C�h&�>������_)���;��i�-�Z�p<���QLRl��ێ�Q�xr�0��`Q�
�]����'1P�=�2��	�_��ĭ|���C�7OG�gI��b^�m���ƚ�h���Ȋ�tu��N��R:?K7�p'�nR��������%c��2([!�u��.�:�N�h��=-���#�Ǽla�.<$��n���;KT����(�򔿷��6HՌ`Ġ�2ؔa�}aM�B{�q)܊q@����FQ�ڨ�o��gt��y�P�$�#�ɾ$0����
�*����H~s 5c���xI��f
��J��͓� "�1{�+�!���|x����@֫����J.�'���@��:��ϙWJ�/��%>�a����jP��Y��z������_d�Xd�5�Mh�Qi��Zz;����>�S����_�d����7��o.kR��ƽM�Q������v�w�O�d?)Կ+�~���P	��P�1���|uM�bG�1��&�ClO�O�ѹT���(��f����kou,ZS��R�>�!۽�	m�CHCzh���B3?[���rJ���-V0M�	���D`$X��c+ l�V���n����l�qi��X���� �F36�Y?�M�hqY��l�L���d���t�?��Г;8ˊ�q_�Xr�0�8��������,�m	>>�K˵��`���x��]�> |�:=i���co%�t�(CK+�j�4�E��
	����Ϋ&AY@pn�NR2�O`n2H�OZ�u
�MYj~Q�wkW�C��w�j(�����s��Vu��g�j��{��ԯoͬ�(���V|��7j�pLf���Pͪ�-���Xx����-ʑ|�O}.4�Q/&�MMr'v�]x�B�p�Ж4���I4S�bU+n��#!0��e|���i���X@�������.�g�2���S�����4_�B�f��ظ(��i���CT���Q�R�vJ�r��x	����(p;��J�z���7���N#�R�	@BC�|�(_؎[62!��6=�?DuL2VB&��?p�5c(�y��=��Щ�1��' <��#A�R��6�j�
�b��!sL��,�ɪ���C&�����ʩ��>P:rU�BB�E�H	'/ت�t���>��*�o���ozvۗ��uBz�p�5���\L���>�uI �y�Z�B�L�~�R[+�t1���	?�� �����R��u�k�v�lq4tX�=Ȍ57�T�j�ή7��HJ�q�N���9��;�'�Wa����\!,���J�����.=��*�:L��84��8�Q��c��'�{�I!�;�va*�S,q���S}�bb�͜�`�Ú󩘅'ڎ���h9��,���#�[��|Z�C��˥D�ۓ�;%&�^���\CG2��!�#t�I~y�ۇ��I�)����O�C�P��u�L�pS����t,�*��­�"�������ۣ�Y�u��oZ|�dw�(���|���h�b�P/4jw��F���� �����}����A7�@n�D�s��'�vD0wU���)q Vn���
5�=��;I����|H�<6v�8S��,���8@�1���̵�n���^��ų MDĸ`U&�'�±t�e�AЕ�'�Y�N�R{���G��EE����8W�<lo�_�F�qR���Ϗ#���b4��c8Ib`�B���U�����2a��A��169���<�6��$��:s�M�?�?�uJ� ;����I�]�n~�/tq��_LW=ÃKp� 9\'� aq�+	*0��ƭ���"]ȫp�J�B�$�i�=^7��ޡ�I�׏t��Kp��S�94A�D�J�,�Zy�Bw�ك���Y�����6�Y�}�6M�Dg��&�(#���Ń@}�Չ��M�CTDx4�)⻔�v��a����FR�1�+D��S�� �~����D�k�ş	�w�J{����%g�N�bSR�[������m��*�3E�*�;q<�q����6|��4�f��D�ӑz<���i�C~a�p&;�{�B���t�G9:n���q�v?��4�6��4Ú�PS�gi�����_�+@�i=�D9��>��P\�h%���.Yc�b�jVƑԚ�` IC{]i�Kῤ<g�p�A��u�0@���x$O��E�L��F�<��M��<�k�]�z2h�z;��O�[���^��~�{�Ͱ��~�����t��S�ź�lq{b��aU����87�����.ȕ\�[w�\� ��Uv�j(zT��&���h���p?�3ȶ�����(?���!�B!7�3��:fo[/�����(��n���S����L�S�Px��[XR����36�����i��(o�`�$�υy 4��jLZ�����PKB���Y��ڍ��,U��3������o1j�bK84qv'Е̿�i��jb��M���5ⱙ&��%���07+0�EfD+D�)���yW��\���D>�`�p>�r�Y��F�j0���Й��L-k���A;SP+�Csf�l��F��_|V��K凉���$�9UYܱ��7#��� g�^Gz��R�~�\IlD����C-O�G����(�%�B�Rc	O3o[�xG��:�1�+��͞�(��c���2A��%�ˈ �h+m؄��=�%`T݇7!��Ғ��:�������D�-MU�<L�u���A��w*�5h��]#�p�]�2X%��~X��)��8C��'���ÎȋĄ���S/7f�Ns�����o�b�ڀ7^�������J)F�nL�9���U+���#:FA�.sF� ��ފ�0β�~GJ*��z�jh�@������N�7p~��>�{�Jwp���3���˃{ra���`R���	5?D�g�ME.�d�Moҧ���Uɘ]dS?jU<��S��YQ��(��h�cn�u�[7D��jg�G���E�9�����������ת�<�/~|��C�P��y8^Y�=Myr�LZ	��ݫ�������V���/��5�N�l���H��@)������"#�o:ˉ��]^�l7�gQ�n5�C%hRmR^˓w�ī��V*�vPW,n��IE�y޵�}��c����P�����Н�"���`��	�3}���OS�������W��nb�{�(���O����y�X�`�F�>a�1�s���|8�gp1Mgb,E��r���틓�v�\P�%�w���U�Y�f@#��������zUD�t���k��4<2!�f��/�b9[�>���-Y*�Ϸ%r���*����}P�4M
�z�����Y���=���t�:ExF)|�Q݈��Օbi���~�e�� /�x-�*�xy�z81wh)�;Oh��|�Q��M�=3��ғn̰`RA�n��`��O�:��13{l��\������J41a��}����?\��]�k�o3~f� ���V< �W�f,�w�G�YT{��h���F�M2��	�p����Y��CO!`����W�kUK��v�Z�����`_(�	�C�����|h@xQ�~�5&�>�t7���N��>�|:1M߶um��06�?�J�O�3 S�M�OaF\S�ic��2�t�ڠ 1F	�*
��EkL�%W�'1�:��[6�����&�L�8�Ԇ0�Ӣ��`[��`��y���=�!��SM��Fv��xqb�S���إ~+�`<��[�|&�]O�N��:���(y�7�V�a���_.����50Ew ���0��|����Ѥ�����n��ڃ5�yK��bf������gUȵBQ�QK'	a!l&�����W1�����\�;Q�B�*=���P���@�6U�ď՜�'����N� ܱNd����"c^�R�EL?!OwR�o���Y�>#�bh�@}Xaؒ}�UX�|]��I��>�f�ᕑ&�We�n�`J^�X��>�N�P�{8�ڰD�_�^�Q<`" ���te�"�� Ai6ﰓ"���J6"JU�t��S;�Ь�o�|���]Q�"NGa�F��pqb ��i�����S0�Dg�I�kP����I��o���
v����w�-�!繖i�y^(�Vc4ʞ8e���ȟd"^]�C>�:׎�/Fp >��sތ�g(vؕ��`Ā�����ȵ�b�i��#�2u�6a�<w,��,�>�����ҥ1	m�[��h�Mp`�>�>��ֹ1v���z 'T[���7ϻ�+1e��nE���j$ �˚ٸ1��<��jDo* �]X[\V�;�"Ō���qi�@�dm�mј>P�b��B�"斮�c��UP�?�A]��(矩Me'��V����e�}��v�1$:v.�P�D0<�@���Ӄ�r��[8���No|��V�c>�oE�0B�����ܧ�-��w�j����<ȺwB������w��������l*����o.gJ�L��V{��n�b�VZ6q�ACj�?[�E��'�����X��ƺ�����Q*��P�J�Р�9��~�!{qX|�O�w\o�I�%݂P���')m���$�K�&1X8L�D%>��M<J�C��^
	��O
b��wiO�%��&�شm�Ė�e��Z�S�ϔ�Z�]��b�fz�w��Zu��c�_҆w���1ԏ���E�:*b*�sR�16v%�@���n��Nlf�N�d���E�����1:�Q�'��݄�J	����Q�Y��iZJ� (��y�����gqĕN���Fj ����s�\��s�v�̥���<��ߌo�|�RD!��w���$� k��P�חYI���k��6,#����݀[�֌��7q\��"}L��w��G�3直��U��a��9��tZ �\kU1��,G7���d������y����ǖ*�����z��"CV䩪h�ǚ]s=?v��V����������s������[�/�1�����̒�G�u�?)��bӕ�/j�q��[.Y]Y�XZ�`;3�ڊ��Ys�7L�m�*�"��ε�|Ĺ+��+δ�(�9��o���>�vfv�X�)|�Vg���� Z�B	Ev����*:qu~y<�T�G��:4�ɀ��z�	��N�ud���g�	&�u�՟^����.�Iud�C� ��G�vD۹X0��s���_���@�;��+|c3�g�Fɿ,`I2Q��&c`a�'����l	#����6��R�7�߿�~��>��f���.����3)�9�Δ���R�����^`.W�������l:��OS\Xg�n��9�k���p��aSD���(�U�Zڟ�ᇾ
>���-,����	�J�(�\`���{Ñ�����p���:9a��n�� L���}������~ �mm��r�iτ�TN~���Mt�4�ݡq*��%����y޷T�٪/�
W%��01k�[�r*����(�1L{|Z������c�[�+�(ܕ��~Fy�X�2����*�i�xڰ�����㋔���t���m _>��	T�f����8����pd���l�)�3W�wH|��~��Ȭw����m�ɫ�%Rgqͦ���4v����x�������w}Gd lT�9/m���nb�/�d8~�����z��o��'�'�>�w�!���7X�q?�j�h�u8���a&��������(T�͝���	m����n!�0�m����[��߮�ֱ�_bާ�td5�Z+ɿm�
b�G�;Sb&��;�v�mf
,R��S�������~"�>�&_�rs|�8s '�λ��(l�8Vu{v�(|L��$i9tO�]�%�Mgx,�X�C�h�ِ�N�{<�ݴ�x��7�7N�<]���>�������d�	0"�d��[�1.	n7v �L�ƃ�-����|���(փ�y�AȨ���}@��8u(-pU�/[��ߧ3T�ao,��$�ͩ��}�FF�����mE엓76(����W���eezR��f�VP?����0�����v�{R��=�N�h��:�eBC����^��֫�$�O�>#&��5��L���>�1ߺ�>gʸf��fa,�5�)/K��Gl׸�e��y�� �1B ���i��~X�"��G;�[�K�j��T��ʗ^�FNi��*Yb��*.v�hYē����gL%,|{��_��t��4$���lp]j��C	��/O�sg̺K���Y�)BC0�<�x�{�A�)<��`e;��B#�Y	R�� �س7|4t��sU"��&})�/z�!�c�y�I`_��1���{��Y����t�:[ܬ�V ��z�w��2��ÇE�Ao+�͞�ƺ����?-l����l�S���»�E��`����� �[������f������X��H��4�3�����٘v��Tƾ�?�,�wf�������D&$�ۗG�ΑL���}��T-�I=ռ������6��4��1��W�M��>���1'x�C�|a��PJ���G�j`,U���`�d�\V(]>��R�L���Q$f*�˪;?'�0@'u�\6��4�c�c��{+����(�2yG���=G1۞���u��Y��خHFx\L�/�b�d�=�G�H�IX�V3OV�u�l��q$p�
�#���Y��5|[�qn���H�X3/��{YO�-���kx~4)T=s		��hٱ^�*,�돓"h�D�xA�Z����+a��Ǒ��{[��9X��P�Vv����<Y�E>�q�,��?%�U?��AL�#���T���B�(� �g9�
s���$�ݲ#樣������7]��pȔ����cU�tgZ���0YW���(#n� �s��葎Wqg{�8`�g�n	o
���u�s��1�9�^�3�1��P�?X9��%O��Y5Ĩ2�Xæ$��A���M΍{�Wܚ�8 =Z�"ߑ?�M	M\��A����
�vWf8��ڂf�pҚ�����������O*Ѷ�い�1Am��jXgu�;���2��KC��_��5�ܐ��\|�v ���eX����Z9�j�lt4�7jn�8"�{�?o�5��D˯��6�e���+d�L*��4������+�|�z@���/Γ�)hC$x���N�l$�uFw�9#Q\OI���oO��>�<~��3��ۨ�wH+w��s�V���wRT�boERo���t*���,�{�=�y�r3T],x��s�oٵ����j'!����M*�~�
J�+�ߺa�?�:�ˑ[.�vO;9R�ܱ!1��h?\��-g��Ybr,��wh��S�����z�ex(:�~�X��Aw�|�x��;�8eM�>P
�f���[������̅��E��4�䡳Ę�:o[��~I'�����G�s���[�� �~B� !hBL�W���7](ى�9��Fٳ�(Y!�F���wq.|��>1�瞄d=M�4s8�9�5eu�rv�/GVh����''�zb����a�}f4��a܃�}Cg:t�nPΉ�D�k�]��X^]���.�>�:��≆{j���߲Fi`LL��u�Vb,i̋���	Ю��*kR����3�ʼ	�Nm��}��ҹ�f�>FB�ˀ|��L+��u�ۀ��?�qm���N{@o��������b���:3��=���_SE�`���%�a�Zcd��t��#R��ły
be����4��)��B�nG�^i���o�����\�-�_�.�j|���`���Yq>���l%2��a�ۃ�Ws�U#ɽ���6	��ۨ�U�;Ҙ�+��Umt����2l�����/���J���gh�98��(8uP����M!���cTO�Gb���`�=Zg�E���Nǚ�׋\[_����#�K�2��^��O0A�~6�S[��2��B����<�{ ������t��z��5�Ndå�1Ѩ� `�m�i���Ds�	S(c�@&2Ko��࿄v�nC����Х�����$ADܺ�>��x6��uh�8E��R�����ۙ7��V]�e���s��m���C.◷h8�'�b�퇀�:NU��슏箟ԭ�#�Ԝ�C�%�z��ͦ��0�2˧�P{U��4L 
�3�bk� �6��W0@��_/맼ݬɀ,�4�?X&$U�#PmmE��,���G�@d��@c7e�ˇ���(
�QF��d��&{Pu�^&=��B-\ͦm0�SUT��Q���i��_U��*��ϵ�O��_+b�D���
�Ht�[�Q3J%�{�~���'��&����L=�9"��	͔d�H8:o�N͞9��C�
���~k}J�y�P�[�Z���J���l�$鸚�U9q�K�,B���?kl!�4'F)хw}ҿt�/��<#mT��a�a�-�LX_�p�X%yn0/����5�^���P2��0��t��2�\�V-4�X���e�WFQ��*5[��d�bɨD��Pb��M�+�#S�{�n�)�V%�̳*s��{����;C��$ȧ�
؅�$��Ƒ�_y�d׼�Vm3��;������	W�Bn��c <�
l-7�P��[�i��1�H���J�s~*��)d^)`���wH[���U��n��6�QF�NѺ4Lk��/��8���ҝ7�^u��\]�(I�R��aB�:ԫ�k�g��b�9�C� ��x�	K�G2 w�<��,��{�s6W�D��o�7.HfX��A�9���7~��AC^UN@�����:.|�GG���EE"�z�y�\�+K )/���`��1(�D(��l��`�t�&n!Y��TJ|�S�`^�Jn��o?����qkU,�v�Hޥ�͌���s�U�[c)TM�t�i�d�����Ꮄ�����ح]]��2^~Ĳ��5�^�ݔ������gp�� U*S�ݖ�E��l:��˛��<�v�&îx��Y��O�p�T���f�Ώ����2-���(��� ���VnŦ>���M샺	��/�t;=f�`/�N��v�hN��|�.��Ǫ��24)�EJrd�H���Vf���z���
�2�[���3�$�y6��$Yp~I��E�����YL/�ⲅ1�v��f���z���h�Hha�"��3�Lԩ|V�RW�z����9�w2!ٸ6B&sa���/��Hi!٦߻UV�4��H�b�|�~��_˯L���zO�F�����Gr��0�!h����gK_��fɌi_���!����c����s|���-̢J���4���T'��.�^�9�qX	��Mw��2M�	�*�D�,E|�罜�swb�C�P��/��Ά)�#t{3`�mdn^������:�A]�</� �S�v7�w��AbO.O�"ͼ�!�l��4�^�w�8�q`�Ȃr���&e�g���4JƟ��r\�'&�qfoሪH�d_�kN�!>��|�JP2��hZk� �C��>Y�i��~�������_2$�3;7��ǎ��ߠ4@�3�>�w%�,:T��U*@����y{M�X��;A�Fg�W��f�6��H��tK�p��tt���;�҂�;�m�����}L%=�
C�?��c��A����3���tTg���\��I�r��|/c-�a؄��H�X���r;�v��f��wQ�K��-�`�6�;�(��CaM�yh�
,S�-�բ��v+��W�,v�3��÷1�Ď��q@�(�n~��c��h��~�"l;Ȥ��S�����\�
��x��4�����H�y�aS@��3A�,�m�"ɒVa�*ߜ
����[W��q���c�H=��0+΢�jE�u,�'Uf���.U^rLf�t��m�J�a�>�FAM�]�����º��u�����٬jFi��c�I-:;�wEg�oZ��%3�5a��/28��0�գ9�ٻr���?e_������\��
]��^0仍�g����^�p7��]�q��~�0��G���R3JG�=�	)�Kc���V�4�Y��k`�o�G>)���j�����_��v��jOҳ�J�j�I�Ƴ���||�P��e	�v�q�|��	�T�Ѯ�H�oxw,��Y:���	6-?���W�.j���]��g����I>��Ή�e�v��ks��c��F�d8D\$�g�n�_qon�;P���cxoQ0�ہ�e(6�R�����=�����J��6��"MN��n{d�〸�}*�ȓ^��E���

�$���\�=���F���~��;���F@|Lu*�7����jfũ���ƃ��3�&*i��@)��(���a�m@b�<���-o�4�[7�?`�^�֌D��&�?�x����_a�@f����I~	���#�����g[9yQw&�Jq�4kBz�G5�Ѿ"�s0M%�t��#��<=k��#��gQ�ס@�pt�ga���k�$��SɍSp؏.>�$�TQ�G�\����O9�etX7���8�5�&7�-e��H�3�����e  8TÊX� �L��u�����6%W��Ii�Xr��j�ƿV�%���K���5����&0Cܺ�6Yb����M�]���$[�/��/�������$Q���sP�\��9�PN��L��-'�s�1��$v�ꌕ���Nǣ��r���7��4��W��Dm�[�q�W&��^o�_� ��ۑ(S�j5��ԍ+�{�Q��E\����3�Թs������gΕ�tP�H��n�,��Af�ե~uɔ۲$͟��p�yT���op9�ly�:�G[���뼄�-���Z�D�I1^��MS�
eٛ��U?�/�t�����4��s���T/d`^4��&��g8���ZD=�.*ߨ/�JaLfu�4�[�ї��)�F�Ζ���6��w�V~z`��k�VB�W�u%iU ˥��D�,����ޠw�v��T�]�2����?o4�Q>C=n6]D�	�����#��/��:��ꫯ�y+N��@u}��&5��v8�Y :0�P��hk���J����MO�t��"$�W	��֦�B���쮙c�iZ���a�J .����<�k�� ��4��5��:nW^�i��'�l���۶�^V�q�>�&"�!���OJ�y�G���L�o[#��[�;>R!N�m���Яuځ]��u_�5}a�~�7r�k��
fzV��u��0���=�K��=ؙ�æ_s��:��t����жH����j�qs1@r��w��#�%Cw�I�~EB3����b��²O!����z����ⷸ�꿑N�O������ZCrf<G���m��@�����Z��DKV|�%�i�gE����߂���ρ����H֭�n����9�k�x+�l �+_R�>�˹�{eD��!��!�vl�TSb��s8����
$�=}��(
�6BO����ϋt(Z�B�sJ]���paP�u\S��
����W�x ��?�_F�7��l�W�v|��s�izSz��s9T�-�_ƍ�e��s_f�D�%��f�hFVV|�0ݜ�S��+vO~N)sMoU1��W�+}j��c�� r����c;(�`q=x��cU�rM�
>/��'�'�4�w�>vԏ�鬌�QZ���a5M��gVx�\:�\��jZVs7Ԉ+�z�5����*�(YZ�h{PɆ>�����MKz�`�		���^	P�^�Zp9��6�9�Ť��~��n�>P��I!����;�������q���4e��x'�kȗ��*�4\�K�c�/� 7�s�y��;�TG<z6Auj8ur�h���១0��Z�6�ܲ��M��fc�	�%��q��̥2��lj`a<�2��u�,� �L���#��E+�(?F�5�>��쌖����Z"����#S<N��2#�i+�x b�FR��Z�F,&&���Q���d[�6������U�t�� ���s|�����j4Xq���k�6��\G�p���ZK�Q@���.
���M���I5�p!�>g�V�l�\�4�d���#:�/�ow�w��KX�n�҇���T99R��u����iSZ�(��2����p8@����=���`��>�Z悐�y�E���:�c��i-�'��+�����G/l�
�{�Ef��L?���B�]��mSY��$�7�eAF|_9����N����c�D�Q�O�(���>�s��s�Y�t��X{E#F��#[��;��=�$wW�/3`d��
c@����VRvb	;{��e�ta�\���AS�SbO�An�����*
8S�u�Hx2�G��$%(�� ��<��c��	"T�'闦�ʕ��pCr}�r�Q���-G�G��՜��pz?��w$�B�)O`Ԫ,�e��#�ebH8%B��j�3`
"8U]�K�z���O$Ź/
�P>��+�ob�U��ւ�t�5���@�+�K��L��AȠ�Y�|��e�����k�v�j6��S�I�������ͺc�]�T��W�p@IZ�5 Y�ȣ#�f���}�w6�Go���0�sZ�M��%�tV�_�p���D�WȜ��Nuk��?+�(MH�^׉|C�!R	��'	�?�7�=��T6&|�a��Ƀ��(;[��T��[;��t-ꭣǵ�  ���ܟd�e�>Sz�-ѕ��ʕ�pyH86��;���.QN���Vm���n��L+�J��C�7=���gZk?�"�u���@�0��3�D.-+|�{�JSN-��F�M"/j@���l�P	�y8��<Z�19����y���T�>u�*lQ�F������<�P.�L %y��5�;�پ�V|H\�Va"�zyf���1�������|O=�^ؠѫ���Y*2YF!6| sJ/lHz:T C�_	�'�h��\M1x��	";3�����&O�7���&m��I��j��!t*�a�
P��~��}7Ǝ/ӫ@f�H�i[�w�#w��h4��Ў���G �oTNs�3�����/~Ղԫ�Y�1-ɨ�.޾{O&=~b�渴�]�B��p�e@bJ6��N�#D��vBY����dH��9�ڳ�6�s-�NGi�)5/�r���&.>�h���,�cm)e����ҳ�8�ť$��
_�T��Z�r�GSY����S�^�=��Cټ݌� �Q�~�B0�4yl'莛E��S���5������:o+K~�)�(�F�8��B�����&��;����W[�2eXl�΋w�-p� ȼ:9�M�Nf��C���kd�0p�����B}{��$L8D�
��q0����<�ѕ&~c�׻��l�b�䠵�^���P� ��1����t��&�Q�zvU�k['b���랞��m"���Nx��l�û�mfB1�vFE4z>��� '�*@p�9���{����01%�dJf3�2�$��B<�2t&�"���������)7�%M` _���lB��)�B�Z�w�4:7)	�[�cL�4���{/�ŨJ�q9�M�p�t1d�`k�J��� �Z�䓹��?���xR���S�dr����=c��˰��Ȯ���C����l�&P�9Pz.��U;���l�A�o���3x�j���9ވ<�.�H�����Cv9B�D�$��L wC�����Zw�����",~xy�!��c���J�+�t��� NDr��ݙ�\K��1�n��L
�(;��E?�N?�$H$���P��g�&q��%�2y�Fܳ�J���@���K[2���������юl�O�zW�먾E���`k,��iS��.�1�c�Yi�&�z�߿��DX
�CV����"�`��A�!PA�3��Dc}�6��ל��'�W�ظ�����;�q����R��ϗ�[D[V��L����0����T��m�.~k�N��GC7R�ç�us�>D]���e�4��ϑY#�+��A�'�J9G�{/o����)d��_����c>�h��G��i�z�H��u���u�Q}�f�U������d�$�Sb����n�V��K<�5��sс��l�縜ȰM bib[$bs��W�����aǐ�E�t�.�|a�<��^_�;)!��&%��z��"�M��z�PV��۹oi��A�,�^c�\j�s�[D��=K�ܻMۺ�t?4��h�̖S�!��KrU>��c.(��q��N��0�*�p�N��n��i��7}�㵼:�%�f���܊f�KB�o�w���qi��^�s�逭��ZÙ�0o%P_�O���B��%n��@�Q�X�7�,��k4]�����tI�zA`BE��5��ľ�١��r�%�_ C��n_��}��D�i�ei�As�w�w���+�x�;Z%X]O@Z��r�����FN*Y�w�i/\a����{��]BUj(��П�����	7$��a�J_�_����Ǣ��;r����1f-��2s�&�FT>LK\�Q�C֎�?R�P'���n�����ن#�:�����y��$sM�e�$?�u>����>��+c\o���6"_�>6t�wf�����
��Az��U�V�@�����d(�*cA���K4�V�.*��Y�<dc�����ɬ���/���^
���6KK�o�r���]�NN�MNRħ��gP��C���+�t/F�����V�X�j]6���yA�?H)�<�0�i�z|�@��eJ.�D�w:������	+�DC�c�k�Oq� C6?���=���<�|��v��Bv�
/���*�v�`�����E:H���tm�Y/r]u�ΞOdI,�8�D�ܺ�\�T��A��jj�/E�Вu�ѾbL���8���i-��a�	z���u��)���>���w�F��ڻ�}��њP��XO�Òv�����L>J��*f��iÚ��[���"��u�bf�RC�2z�r��a��2�'*�"q�U5ort�'S'�E�A@�q���́%�T0�kNi�^�b2��YAJX�ê��~7'�������*���bL���j���-_�b`���Ւ�W�5��T,�������!
�#Ѩ8�6�5��d�k���XtN|,�-*·���;�4s�r��(�rm ��uI��y���S��A�ER�I������J{}v���m��\<`����=?��7y�����g{A�K�r\�=U���B�7PK�%�Mm��p�[_F�,Bp�����
)��Z���y�L�=�ϧ��V(����%����&S="͉HdWN�~s�w�^����9���@��ǋ4�M���uJ��G�UѣF�����w�����7޳� '���P�tzlS�D�?��2�E��̈́P�'A]P��Ck��,���� ��Y��̤̏�1!WG��M2��P�qծ�~�����0!^w�
w�Q��w]ѱ����;���FB�7���e�Sɖ��#?J>�B.��[t�Sʏ����E�ǋ�O+ޫ0Z#b0���%*�MSm��蓕�,��Wo���7<Syύ���r�XJG�������Ϸ�+��A�%M��Ls���`�W9�BTi�b~|�i���H¥�!�+�|�����$�c�&�:(O��V[�6���Gt:�҃ԉk]�䢨f�ķ2#(�Ri��zxT��/�	�e��V
��f�,L prsY����!��p�A��[-�2��)�]����"��_|%�˴�b�O.�z�^*�O��×m� v�Z|h���_��m�&�O{�vq�i,<�݌e����f̭m3�Ë�X�[��ۋG����G覑7� ����
�	z�4>x+�h���Tr�����"��C��|��%�!�k�$�uE��h�x�ԵJ��&~��A���զ���^>��_�{6#���?�u����9�J�0+e!Ry@�D��t�BE�5DcK�V�p;V���kqq+£=����U�ͼ^	��;'��:�'���c� �k�_
h�TG��\$��\V͞Dpl�Ka����y��q�i���X����,9�"I&��Gq����5tw�l�A�E��r�v�y�Z\[�� �<�J&��&>���'t{�O�
غ�t���/����~s M�Z��煖M������S�{�.ϙ��D������h��Y�1Mp���|�ҟ98WM�['�J�����v)':u]�H�j����0��hmJ����౾7<Z����ov�ݸ�cY3���.��d�9c,�!��q�}%u� :G�i���C鷳��;�m0��9m��k��aϸ,X©6;��+���,1l�m �����\+8�͵�Y�[򪐢�m]�VF������(�s�نY��̆�+��V�{�>��s�A������p��zP�|V�'�$0�t���[�L���������NvSR5��y��6@R泷i�{��Zt*Bc��cKA�H�DI�ɟT���+�E�љ��׹!���89K��k4�I)$χ���2��i$���/�d��H��:U1
���i���yoϪ\S\/���3���<�>8���/��C�����>��#�{��A�����"[�y"� %43u
�6�������Ђ�r��":w�t�G��6S�j ��N��8 �ڜ��Ŭ�:��]niR����t�zy#h���Pv�).�5�;���X��?�;��$@�������:���({S��J�An�>�~�O���Qn�	���/ɓ����B�~�nHxL�1@�Hsܛ�C<��<1�z6������愠g���q������ �)s߂; U�R���6*����k���|#�v r��A�kvRJmf�Cp�b����-%�K���E��R�������1��ߺf����RY������G��&B��J'��4Yw�1lc}$G��������X����<��{I�P��J@���:�]�@��~@�I����p	�dph�'q<],Η�M���2.�z�˥_u�9
�e�Go1"E_O�H��FFڹ�r�{����'m�p�k(2���6�<��GN�y�Ω�b��S�,&���q��IU6�ف8���w��l�N3B
�! 3�;RA���
��8=�Q�d���0Wlm�L5��S����
@�5��-�<E��{l���ܛ���!v=V�V��J<e�K�R�Lsޤ�9.<
&U�u����a�
�<5�B�ԟ�5v<M\����٬�
��,L�-xH��-�A��蛃�X�T�7Ѓe.�N�=TJ5w ���	�YfW�X?�c�m��j��Q6��q�x��Ƈ4d���B��8�u�Y���r�3����Ef"�
�p�.�o��!n���e�?;����l�G�ݸ�v@U���/�^�hz�o��h��[f�wڦ� ����a������w�����(�U�U��kF����>z�+E۶���qVͪ_m��'ĵ"��Cy\|�o�0W�̐�^�	�ֿ�'d���	���R��9c4��L F�Ԫ�V�6�ɨ.�������Dg�][�_$�8��
���؇�>�����^�2�sp2'��+E�Ar�QI������2���7�x$
�������Km��NÑ=C;�J���[�V�N�o���iBP~�PZ�r���&�y�)�������t���YA%�&6�2���,�i��<Y�"�=�"���uewF���gC��r}6����|M�TR�s���C����BN�X|��Wٖ�9�VL;e̘�R'F�+���t�*9>B��#@�xU��e���bz4lW
�D�^#oR���.�6�]�l>v��ƈ��`!���"�������HR���\L..:1x\Z���ٹ�:�x9���U����Mt'�0�gV��"�y�KB-!U���,�#�FJ��`��� �VY;,	��B`�%��@SB�"��̡G�y�v����|��G�g[�;�Q�sYl+�9��@ob�W��4{BS�T=��;��0�(���L�˵T�Rw�\�5�6�g耂i�׹�fe(�h�Dd;����`�&����%�gi8>���`�:����}�������𰐭ܵ�b/��xN:A�	�ʕCJ	>�V�8�9#�����~A��a�H� ^�����ɛ����:����%��ֱ���4:�~jЉ���)+Ϫ�&�A�q��Cb>�7W���IP�QK�o�����y-��:�$^NkLSRT#?�����X��{RG|��L��r)V�#oTWL�v-�9��7�ٙ�.f�b���C��7���z��Y�)�=Bu���"C�i�Z粠������z�[�=\-��]�b1�J	�Z�tk�֌�P��f�r�q��^����C�v�aX�H�Lx����uVbZ�9���D��x �*���?@�XB�9ү�hǸ�]�gEԘmH3;�O��z����3�c$|/��塀�.�`G1�8~I<�z�DYQ7��&l�����eWs���A=y.�Tp�p���{D��e�$k�{( /)楸~�j�m%B�b8MP!�ۅ@͂K�y�q�8���d�[�.��"K����q 	��K��z����5�H���h�*��5v`W��)gr����`��[y�Jo��x�G��5�8�r/h���'���/���O�QO���LN^�k��F�s5^��M�����Bx���ҼL:��"܄��!�@�]l©�H \�sn&V�
|C�xѥ x4��([Q�Y�bc ����l��u��1�_&��� ���T�Kb���JW��'y�$E�&��O��$%7�ѺL/Y]Ze�&��&���k�WWQ����s��IXm贔i�L��B�T�e`�o�[iV��q��vh����/�R=-+OhVm��ۄ��Qs~�ț��&��+�F���xF)b�������?���\O��2=�3M �m��FD�O�����̅�����M#_����c��(�u���xC�$�&�Y��+c
��$CTJ�u&U�����'-S�:��>��K�u�<�Vw������!����x�*�A5�V�b�|���$�&]�Y
��X�kî^ܧ[�H�Q��Z9!m!��m!9�v�^�$�o����s^����i�
y�K5�����bY:��Ei�x��&c)n������̫C����8�L 8E+`�nd��%1P�'�o��&�g"�WJi,?��:[֝�}�uF�o��KD�#M�����c���_��sЦ��m��j�q���34���U�a��@9F~�|��Ȧ��\U��gE��$Z��On��< %펁�����I�Z/��V��=�$M20ܽ����u��N.�@�����y�'�Ա���s&L�?~9?��؆ .�S�H�u�`���[�3nP�f�SsJQ�oԓ�����[AH�y���2$|����,z��j��[�^�X˷Y[�A~��T��ܽ?�U812&{��	z��>�eg�	oO4�ϱ����x���h���t6@�E���0vX'�ϑ�\�uw�$;��z�r��ѠF.o]H2�L���\�0n�P�)���A��+��e�Y�ٮ�܈1.<H[Щ:�/�"�$/H���/F�H#�	�����e�;�cV�CX�O�Za��i��><�ZP�IN����]�Sz����c�����$$�/�Wnk�����9z��{���pߡ�/����WzZ����I��8��
p<��� �ϫ��	�<�*�$;���m#�oX�z�M�[mv���;#��)����LBӻD��D��J�>T�F1"���9��~�ά��}��G
s8[��7�=�r��o�p���ډ��	ݴE���^>zRb���!��C�J�W�x}Z0k�h�D�D�����:�=�m�����C�f��DȻ�y�X�J2��Px�{�C�	U'@��wB�9�ze߲v/��W0I�-��C��"�����/?ETl���0q�%ͧ(�P�,Fg�j��ȇAսK�˻�6�[X��P3�ð���ncн�)
�$��l�?	�`�'��o�|Ɓ#YO���To-y.	��R^�^��[�ʽnͨs��Ld���@��r�e�Bk�nR���FW��q��H��W�/��x�Lz�/t�� !��߶��
�<���&0;�.y~�'	��m�W���P��K���M4&�1�`H�����S$"ʄ�=�7ڈ�B28��Bg�|����2����mO��V)	�B�aY�����3_0J�i��%4P�?��ލ��I�t6p8]�<=�4r-�J�j��Y�d���P�o_x��u�'�N�:���I��52����4���F;�fxKi�60�f��n�������|�F��]��1���ҿ�Ā��6��
&�/+����*�Em�Nn���]�KM|P�8s�y�T^���C`/�bE!~(�$��>�vΐ{����ҶW�F9Q�N��xV{��e���!y�B�����EQx�(���!Ff�߻Zv޿h��W�!�qQXX�<pv�AhH�R�Ӏ��5�����q3d�	�&c����N�������H'�uK�ժ2��,�w�����n�� 2�Ğ@8ھD6��,Ow��p�ܧ�������8]:���{1)+�W�c�n�z�ȼ}�Ǖ\�K���Kz_�\�=��
׷�*r7[��T�,ԧ{Lk��Om���|u�۰x�\�V����{$���"�2rZA���v���X�D���2в<-��I�ɚ�����`��`��%�M���=�!�%m�<~oύ�1�x5Dù`g2��h�.�:~c�g���'��b$��UaٱD�J�0.���Z+�8����J�a�V���l�}3�����s_��~������)ڏf���M�p�x{��;S�T(v���O؊x�3�}kLj��B�`H�y�;^�)1lg�Dt�k�+ �̻]����z's�v�@�G��s��\거�`��
FmZ��S��/��=�,��� ���[�Y�!(|4��\j3}ֶ���7Ӿe_��? �÷-7WxG�yΠ�A{C��پ��Zʾ�b� �������o��ޛ*8��ɭ{^�_H@PYM-���ք+����"zC/��ʾU҄�uO�+�̿�)�	�k �b�fk6xj�*��l��ev�
����+���ܔKku��U����9���}�� ����#���s<�~6�"wc1��:B�h =���0��C_�軽n��!-��ֽF�G���\S�3�f���0d�2Pw�_�;^q{�V�ت�浽�Ƿ)���[^��<�����]La����	��� �R;�4@�3!�3_�>u���Or"�/�iWf3��|<!@	��9�⬽����+Y�{p�Gb���%l�!��4[�4�N��}���O
(�oy&�:��%��P�t#	W	t��/9a�*�X�5�	!�/��BxL�i���A��5�������%���L1e��0"��_I�es��h�K˾]�'���8*��67"BE��0��<���%�A.z�}3��V��#Ť�i����|�L<�dϝ��9t6�HM�&�LzԒwI�0�5Y}�>��ܪ��W�1cM�7��P�����L~N�!>ӫC����.s��?�y��5�<�Q��U��F�d����I��8�*㉲�D����2�f�$�`]�,Y	7ϸ�7Qv������	j�$/����<�X$�͹��*�x�����g�X�g�����
�t\nve������+\B��ԊE����/��i��=Q+Z5=b��UWC;F����;2[�^/<�mC
Y˪zt���Y��4Qx�N�aQ���6�"6sO��[��3��Pێ�_�3��/�I��_��g5m�~1��P�B��.��Ǻ։�ְ#�~�?�ƅ$���[���A�{�f�	��E��3�?�(8�_W�a&QL��%�ې�y���2Z�A���y=J_�R�Ah۶��J4����N�� ���E%��Cޑ��?�fuc��c9�)�g���y��<�[Ć5.�"��os�쀭�[�
h����"��}��_�X?��!|E��C�y}��Ҭ���(g�p�O���#��yCba
U�UqͲ�e�������K�A��lݾZ4��נ�D������HaUB��g�Oυ������>��GFꖻ�����km!�1�j�U}J~�����%���.ӗ��Sg>�?�q��4�v���f^#"��*��`U1��5:�m�`�C�R'��!c6m��Eh4vv�kg=ӑ~��F�K5 ���{��W�C�����u�P��D�2�%b��B<Q�h"��4����W�d�Cq�'^/��C��Ku����t0�	�w򝒇-nq9��k�hg Tk�QKq�+���f�g}�|�\��v"'��S��,���y5���1Q�V���mӳ����uf�T$٬�I��)5�	"�vi)�tɃć?�/Z,*��$y�� �,�g�s�����qKcW��׋��4�î:�˪|^;7����bP�O$�c�<�J9+�cή|�n3o�FM����rod׃U�A��2̹:
��&�菓�@�U��8RRڸ�ˍ���ܒ�4�gQ�/;d�����⍟w ����\���|X��s�[CeI���M2�|f���?�wچČ��]|Ra�:KK��s������M�����m��>ZBs*�-M��ŵ���������ǆ�*�@E���U�A�ɪf�Q\�U�(�5V`��X�����kA����������l[jCx#C��.��2�=����mJ�?���2ƽ�E�[F�%�d����]ŋ���k���sl�~rO��n�!��n��Ӛ�U{��W�8��`A�������?�7���Zy�_�ʏ��^�/p	�G]�C�5���v����[߀�p�G�m�3�WB�6O����)��6����z>
�/��\F=A�ջ�0DW�	�����Z`� _&y��a��j�I�������i����i�p��M����^�TCOp<�XF3wp
VZ��:���Ss��H*�
Sz҉vmv=���6bA<����� ƫ4ҝI.�*%wj��یs��#x�����Cp�ɨ�N{9�`�"�Dm`j}�İ�ACj���Jüwmҩ�&\���m��1
s����WR�H3]G�rd"�;'5?Q��V���ב<�gdp"@�!��B��H�l�'�%U
��Tii��$��z��x�g�6��TZ8�AڽZ�`~�F�8!�嘲���W0���� ���y���x]%ث�h!&ڱ�}�'��g(vp�ZYƙW�2E��ǁ`���q���U!Q-��ɰ��8D�����\=qN��l�A]N��\b${�	w+U���H�rפ\�VϳY\x9��4X�?}
+�����O��rőB���T��sy�b@?�5�׫��I�p*��+<r�����X�:vd7���Ӽ�+�>#ZNL:�{��l�R�^dC1�[�:)9/ˊh��Zg�ϰ�~%�"ι��H����a�_���&z|�2�ꊻ#r*��6V������ӱ���|@Qc��fH".��:{k8���PL�;@Ox �l`W��4�n�=�`��,+@)�3ic7�bgE���Q��K���4 .�:��V��I�X��^Q�]�A�Yǉ��1��`�D���^n�N�u�h��[������`��讁?�pk�'�i����#���Nf�T��F���:߮�i��|��2�b�'�����Q��Bt@K}CbF"8v0��)�x��R7�+6j؆MX �l:-ڙ��m��ɮ	4���\��UnK�Mw���>#�0�H�f�G�*�콹0,���(�	�G�ǩV����M6�ᯂ�ո��'���ϧ����7<�3���sT�T�LY�p7���K�BՖr���X��h:�K� �^��A�B�\���vn*�ǯ�K�9���� ��9!Q�ދ�'~���[��Ol��}���M�3�c�������0FCC>T؋GǷlt�I1<|?�0�\���װf𑣯0C�^!o-H������f������-m5!Hj�ݛ�wyKcr4�Dn���[F\��5�#�=��k�B�"��/�����	�+DF(���8ƕ��H�$�����N�3���y�/k�+;���2J��}��&+x�h��Î�?su6��G�	�&R��V�wl0��]M��E�"Z�u��Rd�"��l�Tp��d,S�l��:�J�(T�>�c�օR$�<�t�'RVR_J[4�~����^X�x1G������5}XJ$���������/*ײ<<�UUM$�i��{.0t�m#��N�ل�[rT~#!mbsX#p���3�`|c�5k`C���?q�zy^\+H:��x�;T�^<x��>�Sfq��q�1bA��.�S��[:�YE0�}@��������2�R�d3���yQ�0�ξo�G1H�7�Ҽ4V�`���1�az�L����?[)	�հ5b^E��7y�۰?�R3y`����0	vN���n�.��:y��JE�F��źoBp�wtt�sk�{�:�[��Ƽ6- �
�h�V�4�1��O�ړ$qF�z1]L�s�n"��)������>w~�.�`c������Y�s�B�$e�W�P�6$N9Ph���5���r��E��b��)Im�@�vC=LT(�s����F�	����Gy�Cؼ�Hj`B~�����+����OXu�(5Z_��N]�zʈ�:�@7G�PX���e�REZg��q�!���H���V�yGJ�
��A� d��PVU8�o������#�e[ߒ5��qm	��N8Zؤ���iR�PF�	�Q,����Q �VQ�p�o�D����p��� ����n����1"ue��X��D�B�ϯݞ�4k����S;�'�"�%�
�&�	)Y��'��*��*F-4���ٺ�{������ظV���5V��2Z�������"v`�L�t�x��/����C��Kˢ�ִs�Np�8U�.��>�n&�zIu�#Y�m��Hn�Ikpw��h�A	2�6�XvA��U3��=,�&%]1<�l�xc}��! Ǎ<�|S1�O��g���+_��w�\{9�f�x���D[��8�z_=�5�(?��Ǵ��u���ag 9��m[�ì8����u��a��+߹��r� ���+��[�1�(F[�D��)�<O\U�z<���Լ����j];Q�������pz~10p"��bqבٔp-Ӕ%�X�3�0L'5v�|;�'U-eR�[bi!��ox� ��sƗn!�Z����7	nKUh=�Ya�/�js��k��3�,�wX���R�f����H�ex�V͸�4�6�W'_��xP�EV�<Y:9������C�>��s��t*�]]�Vs푬VJ�CĄ��57�V�|��Dw�����&M#3�8��r��3�B&?���[��'���S2Sz��`�4�̢�����%�Lb��|�v
�A��(B܈��I>_{Me��$=�Jw�`���W�Zvl9���T��H��d�@�L¸�������=���DwK�.�,V~+?�05�~�LJTt�ĝ��t�]q�U݉�)��ʑv�J��#�y@g�]�f*��I|!��r��] ����Y鲨��8_��J��<����s)�y3�h٦��h`��H&�����"H�f�����B�Le� �w?&ִ(�qY�K�ҍQ����Jê�OI�VM����=�%���5����o�AtG�|�`��v;��Ĭto�t���e<Q�nޓS��W�>^��u�s�IC������Qxh�:�I:&��C���l���S��y�y��rư���6Y�Ԯ��$���7������ ��1'ʄ���\�Y6Gf�nW/@�
��tc2AY[���o<��k�J¹�ps��+�Q3Wσ�(�����"���f�H���R���1���	w-۫{$�va�"�Ÿ���t�ho�/q��|�J�ާf�r��cKP�	��K,µ���}]��L�f��^��a��JG��� ��@�����%p$�2'Z�mD����w5��[��'��cԜ� ��@�����ٓ�=oV=�A��d@K])�^�������he\O7أ�	u�u��c:�޺QA�_�`�:P���	vא��Rʁ��G�gkPi� L�t��lp`�$@䏎�i�=�6�$UQp�_ߝ����G���F�ͩ��
A��v<=�?�}���X6*!��)���ϫ��>��� y,$O����Ō����lȔk�C5<�?�*�eWө˖H_���f.��J�$�໖�;� d�:��r������� MV;X �b� �}{���`���%�d���gӋF>ᬚ�g�G+���]i Y#���36�ۼ]��@��a�i�F�n����ۙ�P�0�rGV��/�u���z�ޛ��X����X��I�$�[E$�Ì���b��
챐}�Vr&ȾKܥ�z!��K+{�1�A��#�I3��E�V2�ԹM	87>��S�Wr3nh�r }�t�q�[O�y��S�k-������C U@�g�SbGI�Q�(*?��;H�7��;;��%\�<黁8֯t��jҖ���G�K��:33#�s�R�BFL(ҡH_��8���b'�a�~=%X�ӊID)x1�Q��=�2�T9'ge�70���z��{�=�^��Ԯ��|t� 8��M|2m� zF��Nn������bٹ�Z����~3�%׌��l�I�����&�������M�UH�?��v�|$��)֠(Ep����:��ܺ�ܒ$:\j<-�#v���F���f$�)#��]8׽���B�xELc,}|���K<��"4V�&��w�6'�)�W� ����t��G���O�H�W�l	o�t�xt��}�vF�]�=��^��S�8�>�
f�n����;N�Yƅ4��b��׷���3�lb-e�Z3D�Ч�V�M�Ả�1�Z\��}y�{�f$���8-�L�L�$\R�sk�ؿ5@�R�C��N�����jV��~�Nb,�l�ZP]��s`u�?)�����jƔ$��kj�P�?w8��7�A�374e���\ot��.�����I�?�U`��=���gL?�:�������ɠ]h#��vA�b.���X��@��!���K���#���"��k��?h��!g~El���7���z�g�;�)�ކ�����wD�	�IO�3�u��:��pqo�\�ޖ�\``O�H��G�gg�7��|Ӭ�Ya��=����ge�>��/45v
T�sA�ڶf��͵R&�)�L���I����9�4m`
�C����~�6��z������ɠ	w��Ѧ���}?Z��(4,���@*�:��£�K"QFO��	��ę.��}�l�Y�x�.sztc��j�vc����F#�}k�e�����^Ud�y+Z�/<��h<C��0T�!Ͻ��r��-�q2[��|%dvG���z��o���X�bm���	�vUc����l����}�1��9��J4�Ǹ��N�';uj�4_y��8E�N����H�u�V�1�9h�S36������re�_��/�����Ҋ��dT�蓯%����RYC}]h�B]�� �-D�E��<��_y��.дu���Ś��Uf풝����R<�Ȭ��4C�D8;ަ)�;�T{���P,�T�<����?f� O���C��)��PMڻ�����O�[�,>_�4(#��w�4��v3�"DZ��Gѣ��_��![&l��׭�e&ň�l�9k�S�*�=�Lkb.��%ܙ #��w�\�����&�q��a�"��h�7@Ī��>a������lp����i������ݕQ2fE%/���5h�6�CX�+��|w��%u7~Ն7g��C^�@{��LD���o�G�Y=ϊs���v+,�2�׮����`/☪�>�b8�qS[�%�Z�T�]�nçJ����/h!U��ۀ��ԩ�Pw�@��W4Z��_�ɳ���_k�x`t55tD�솧�#��^]�� �W���H͖�q�4Dʓ�ʛ>�V�*������
�)dD�hV�����������Q�B[RS�����r��A���Vapӌ%���Cr��&�y��J~��Ϝ��y�O#nF�e�����-j{r�NQ��{1����BWH�T?�.����"5�+ۚ��_Nx}�I�h�=�/JYa�XUQ��� 5`��Y���D����y�oo�<5ʜ��΍MΟDl܎i�^G�x#{>�"�U��m���~SJ�qs�Ō��L���������QL6�	����	y�D�����:=K7�1��bQ�*T|�F����R��`���;��"hk�+��er�'%�!�S�����r��毧�~Ј��)�G]5���X&�\ Mx��"�eh2�1`��i�b��OeFá�c_Q2��� ~i�="@�DiY{n���+(�Q�Mn��7̞�� 	b-�P���1^W��Z:?.��C�ve�kR�@x�jOR���F���V�g�cV��cS��S���9G�~���TH���NÒ���3��J�۳I���e"��"�Gp,��2�9��*����Z�!�&	��=wT�E�_V+gi��Zȷ�4����R:\�1j�g�#G ���@�z]Md&q�m	��;��t��횭F�v�{��n���;0O<M�&5�*}��.���҃�{���G�D@�EMi[2��d`���)ܪHޠ�q�0E���X���6���  OMB��Xj#0�_�Lro��D+V��O�`Q��<�׬	d8��\�/}<����M,[,U	�P �yT���uIWSiFjw��f�����ш��$[���Ji��o��|�`v�,v���=�8��v.rF����ݏ�0��.����hI\�$�s5Njc� ������'E� N~�9L�
@	ݕ��]:lͻ�&�<�#��"���Yg�1�i���Q0�x����VDx�K�@��z��a����"a�O��4M� �'��b����aԮv��L��.�2=�<'/^���9H���z���5�4�5�(��p��,��9�pp�.d]�\rP�T��K^�eJ�җeޏ꣕t�V-G,��˿�!�]#��]�Ub>pS�s3��I3���u�Y*qn|	Gr*=�g���< i֏��Ç�z����JdHV0��u�B4	��珆�q�	�~*��)�w�aW�g�WK��-./���g(żeVvI���u0�2�\q���-�hW�snh�)Ǳ�/o�&Y�=�%��W-�L&��%��
+d�T܎m����U�r}�]��������*U)�DRٯ�DCIc�b�U�z$BM��r��]Hy��5!*H�-�+,2CS�"��U���0����(�9ǧ0�H��m8!��j���Q%���^�w����baZU�N῎@�m)��R|��*���D��ƾ6���{�T��ud�|j.dY�[U�p��5:����btĘk���_�o
T��r�^����+�9��e�Xv	�e�g<u��X�'�*M���t[<&E��
�O%T`� ��з�b��6�P,�_-m<��~g�%D�8���񬊹#(�c���K{����ͧ�ܸ���!yW��+g����� � ����f�\s"㵜�l����F&_��bЂw����N%��n���B���N�M�c;�@	qF��/��v�o=�wK��k?�<��x���<r�0h�[C�J���P����]����F�U&G�o��1��*�#<��k�6�T�-��FҡJ���,p���Ws8�����»0"��2k߼yd$��� 2R�wy��P��~ľx�&5{��w�J`�m�ߑoTZ�K��0}��A
�+`�Ғ�5�L@,�u�v�<+&aR�R���zG\����qE0|j�,t��������EӋ��X�&Y�u���I։�hӌ:�}�++�����q��SG5��¸�]Vg���+L=�9�'���6��Ə����$��Q�?qkء' x�I|U�ɩ�w4c�2�U\���O`#���%$�#�F`�_�p��s��b���� %:X7�r�^ꊹb�q��(XԽ
R�M��9E2Us�Q(b�شF�(���X�Ԇ�&�,�@fS���L���&[���*L��{����4[��9E�c'�*"]���WƝ?���+ �����ݞJ/'	�s�
�8=�����r<8 �k�w:�?��`1��co ��(Y�#u�c(�L��N�������4dV�X�
��g�<q�?��x���
;�T\/�?�����(8zp���cs��궃�ݭ⦄�Cŏ-X��);T�`>�;y���-��'%�u<`N�SDE�P����!�$��!���?τ���-o�Y?&�7�����8T�JIp���j�."�G�T�2ȁm�x_őn��V�7`m�a)��F=���k��#�je3r��0�Eo�e�	|NQ���P[�Y֖��>crwh�vN�$G�������Q��I�%�B�wID��AK��I��'�iw�\�|�s`�]Tc�>�/����z7���`��Jթ.3M̻��� ��;u��S �����d�\JTEO.�w>U�u�d��x�:b���-d"��@\YGq�җ�M%Br��s��=¼��6�)>�����am��dڷ����oY�����p>�X��͠ɀ<F��cN�D� �;���H�_�H@׵@U�,}�J�=Ew5n6�c�Z�B������[H�d�[W���'v��`+{k-�p��A��j^�K�i�5���ë;!�	?*�#I�0A��b�t�D�O��l�^��o��� #L�u
|88�|c��T?I�~�!�������fŚ�A����q�z��s�7�v�Z���X4N"	� 8��[��k���8��#����>�a%�g�9M2�C�X ��`�aEs�w&`��F.�;���5���>_�&]��:�,��\��jZ�O�;W��A�N��B#��������ˀ�<P'}pg6?��,�|��vl)G���+Y(p��&<�i�����qhb!��R�����U����R�����k}�Ս�>�W����o�rz�Iy�	�m�����i�Y�A0(�_����75�Hq�$�K�-p"E�|���;*ͱ'�Ą�7^k�}A#fɆ�6`]A�Zs^}�j�u~W��+ ��͕��M������gd����r��I�~�X���C(�Dn����TǮ9l�o�E��*�7R�;�,�0��Vy%�!Z��~ݥ�_�=��Tf����2%>p_e�}�i=�A`��v�I�WT� �+�����qe��{!�沧;��n�d�d&</�y�nۀg�( ��6�=�'�@0��؉�g���{փl���<c�Es�����~�ɿ�"#�q����{j��.)i�Lk�x�i���#O>&�s�e����]�p����m�3���`E�b��1ii���G`1H��E7�|Ħ�j�m�"����y}*?/���D4(*�������f+ل�u;��\����d,�����n [0�I#t�d`�gc���P�~���P��<�����y�kc
�r<RZ��{/��o?;	�d��1;�[9ǃ��͠�#�f]ɒp}����8'�ۭ^���h
*O���۶~��Y^�����B",�m��s{��Dk)X3�z_�Z+��~�3L�e4�x��#0�r��IE??Ld8?��b�y�'�����*$��ԸfNV�RG?ɺ��{�@���&�6��"�|�`KP�D�y%mI/���fyI�|��~0�:���ϴR(�ﭯ	:���,4��pP��y)V��h"������©F�Y�n9r���(����:��-<�b�$~�����^�x�ۍZUo�f(P�Q�I#'o\ ���&�6*_��t�� ���:�3t��p�Y�ϯ�7.'��;Ƴ�D��$�)�j�)����8f1�
_���FQ��Og�����/=���T7Ŝ� �1O��K�K]�ft��^�X2d9hJ�Fv�i�ֳ��m�M[�	߬7	��YXA�ID��%���d��8�)G�m����J}�Ιb�s�̃X�ā)5-Ƈ�R<"��|,�vF/��nQ0S���+f�:���0��;Z�%8�u�ɉ��«��F��񩞔�I,X3�H��H��$���)��}�Z����w`�&XA�$�O[Nh2�94��qx��G�wS���h��m��`��qC� q�L�~��b��i�_w���/e��3��Ը��f�AhM|	���`?>8�M:��ɳN6�E��X' /S`#�]�9C��aբ<�l�-��ۅ��@7��!q�����L�ϙ�[4��wh3�uK9�+(����V��D����Fy2�x��F����j��L��ẙq�@���$�p�iP��2:>]��l��ˬC���L�/?f���I�}d��
:7�ӈ��Db�C�Xx���#��d��.C���NΔ҃b��ܐE����ܚ'����.R�.xfu�E�RByJ!�p2�z�|�/������,M�]qe�ذ�z��c�]Ù���A?�y�X��u/�0��5o~�_�e܌�;�l/?k�x���Ϸ�^�G�L�^<*Lq��M�&M��{q�Կ��)B?��`s="��t)����Bf�D#م[�;aeN$�ir��F~����vd8r'��=AC�gP���s�/����#z$�NrvY���x��3`��$��e�` u��-:���1I1`��a��Ӥ�_�y�S���ܞ���Q�Bv��Zgo6��Ϙ��L����ɚm�ȫ���d�z��]l�jf������c/]�ӧc�FV��7x�����*�3���$0B�?
��m��/�˺�}�(_�:\Č'7NMתrT���-I8��tT����?�c!= *�����c�烞ŏc�$ ��\W�ې[�ݢYl��I��IW�Gl���\k>����!~�����
��r����U �fN��ipN7?����˒��u~�1WI�l�j�*e���LV��`"���� )��#A��e�o���T�HHr[��9��sg|5�G۷_V�>�lʮcw���ai�p<-5�gP��W]��X۪sNI1/D`�I��1�3���R�,�R��)�n����
O�G?��@eZ�^|�x��T����%��2H��pez��]�a�n�g�֠ "=g���Z����}k=R�, �J!�*���&��yl�*���S��E�g��`�� b�J+�z��B�"-m��h�20�'����C�\���$ B9ku��~U�u-NT��#�.~�k!�<兇�����eI�wŋ-9]n$S>��lc�xFm+����C"t���1�f���Zv���O=tz7h>܇����&hL���,n�&�b��Q�>gmC
�J�~���gJkh�/�Ǽ�ƀ�vQuQ:�B|�_�O�� �n%C̮��^�Nv�Zc�u,B�]D��tOZ��u�;[���?����W�$3!�밢)�[MG������8���:���w�U�*}%�b=�:�~�pw^F"q8sp��y���KD?3.U�5cb���
k�@��Z@Nc�V���X��*��{#�~(�C���d�)5��H�[���̝Q9��$N�O�Md$�V��`�׿B�x�/��j��A���H��z_0��yJ�-�2���A��z/I��R��AA>�����`��N�E��c��_�(�����(0T���w����ȩo��K�*���i)��u=�nH�+��~lv���-�m�����^0�I~kx�ޱ~�8}#����9��ae��R���,���]�f�WZѤ�]8�rg�eki��Y�� �t�&��H��C�uz���y8\^Bۥ��t���3� 0U�?+�ꗼ,r�*�=�Gu�n�k�*�B��wh� �Du����M�����8�oab|84�ߟmm��FA��NhQ����`\W�-�|�
�����ץ�B)�m܉�$�hgj3��9!�<��G��kL!c��)���(*I�V�O�j�@Ĥ��[{��j�����[`�X��8�ޤ�ҿ<�����Z�����Ș��|�6L�H	�ra�9���R�^q���-�$��;g[�9Q�: �G�����N����B{,���~5;�U�w���旳}�)θ�O��J�SyƬQ+�!;8�S�}�!�#��1͊��T��Y��ǵ��<�
�ې��G��EՑ�YW�s�fꧪ[�Y�Z�J�w#xO�N�`�E��Y�&�2���,����4~ꎡ���s"1_�$������#W�݄�[�ۗ��)�������~�È�������ɢ��L�HȆ����w޻��J� "n�|��o� ��<U2�{�P���XHx�U�U��;ǩ���I��l��A=2�A6����I�n����F�W�m#ϭA���S��gȷ�j7')-�8��>�{0%|R+g��
�����^�)���+���g����/P"{O5�"�T�5�����ai����h���)��'�h�1YG�~	���L{n��d����$b�}���R��H��f�/G��е�Y�V��t]K7��o��^�9=����㌖qT���V�������H5XN��*L�*1�3J&#�����Je��z���������b�L�x�y���9��y!y��(�yo��t��ob�	�5{4D��k[,�G�
�����Լ����}pem=�+�w���:�W	��'��gà'
���(<s���	��l4<����j>wD��4uF���bJ�F�H��m��{>���T[8TV���[�=���EF9+ۼidw��mΖ�A�O*Z������X�c�`��<^��TR�
`��_�N�8O�Z��~�s��4oBa�<W'�,��uU{���40�}Zo��Å7�E��O�+ѕ��8��t����̄D���x�RH����m�<v|���|��������ˏ˥��,��gu��]�<aIq���mF�w���p*���r�sz�5���I�G�]~ M��5Q�ڽp3��h�^JNڡ�( Q�4�n*2�{0��IL'��z��o�In77�e�F�pm�O14I�� ������I���H���0��Q=�(��|�80�H�V�"ݺ��!G����mLM>5��J-.>Aw�uf���)����h<�{��j27E�灗A		%�4!���7xu��
U������T6T:�I  AU��=��	��G�>S�%p��W�Ͽ���FT+^���{a~<"Q:v��&&0�%���2�HIG龂��ncQM˴Z����M�3�i{u��*e�M�cV!�ҘiEy X�V| �1��*k~��s�@UBڛ�`_t�����.��[��� �i�r�TΚ&���l�ȫR�Ύ���:��aa�CҪb2�R��@5q<��t9��Bo&�`ϪZ�x�eW����٧��L��U5�C�y� �F�G��" �Ć��z��D��3�-��Q�_�
���IϐO
#��D2�i��S��:�T�,����u���0�1o��t�%�bo��,j�n�FJs`��}��u�$m���}#c����?�>j�~�\�8�L�<��{�9ݨ'�eWDص`p���� $k�M���
i^y�s�G�V���n��E��\�&x�Dx�T����e����^�.fnU��q��A�'�\�WA�B���w����j|���>�� [��#���yB�#�)�p��|(�G
�!��_�Mo*� `���V����M���	g�C�u|+���\h�������b-�����l �_����@u�����^F6�7j. �Z2�s���xD3����𕣿z58fJ��@�Ks�I��n�b�e+���$���|�0��jl�;���6q�S�h��P����dy�h�9���ӆK��/����p{W����>s���a3q����
�t<p@҃�A�dp�ɏ�����L�����
��r�?9ih��3I8d]˄٬��T��fsշߒ�v�$�at����7R{s5��o�OXؔ�K��tCj��<�zJw46/�a`��#\&'c�NIpm��h�uo����l�6N����Y��2J󪂸���Y��X�XLN��a#�Hz0���spg��	�o��*�h3�2�]��Z>���W�)���}��8%*�?�	��7��7�D׾�x�|k���1
��(�s������9�tz
[��w6�s.*'�]fi�e�T�5�w�P��=Ξ��?�f���v�����%�i�Ⱝ��CD�c�q����B���"�.k�C����!
}���8o�(]�� @ٹKv{|�=��W�?��T�0�K�5�D��qI�Z���Bx�Tq�=���G�2�I��:��0l$.��$;���.��אh����9�
:^ �)c
n2$����ިA�K�k���2�M���k��{I�&�� M��&�暬r��"2J� +��E�D��p���w[�4ս�׺Z�z�o 2y���u�s�ř��q��"J� ���VJ�*�Q��ڴh�fξa�	y����i�M�+�?�V��haBK*���uݕ�7C�� �Omn���Q�HWz��8��g�n����V&�|D')�\�t�͞G��;Ա(Jܪ��%tT�xl�dw�%B�c��PC⁨��v�l��ա9qC|�c4��n��.��	P�����e#�G=
����Ԯ���t�8�5	S�D��x�b�4[�L�/ G��*��8�q�"g+����'Dʐ��[����S8B!���<b�N��_�,��@ו�[$U]�4� ����h���'ŉk���A+=X�c72���pXTs����|{�^����������#,1�ۯh��Ϗ��Ӟ��i]BîL=R��z�S{T=2s�=&�W��q��4�Cnv�U��1���꛽����p>!��Nn�F+�7���e/�k�~7Օ���3���Z@���˷��T6�f,^�ݛȝ���A�[��T5b�������2F����[GE�+-�k��Y�S+-�fCM-�U�~f�0�rwa��24�TsC?~?dr���l����
}��������b�ƮA���:�Lk>R�q���Y�*&vf��h�6�5#�i�W��fv�q�f�;l	������4�}��3��x1ɘ����t,�!�s��T���Ͻ'u�5fTzO�He�YY��%`wU��V��	�E�l� �m�ǃ���lp�� !�Ŕ�î'G����͇\���
�i'��PJQ���Q���*9���a��?���9��䝄!v�P�<�t�k��.�e5����)����]�Os�4,D��,���R[hބ�Yz�#�ת�UO}�2��yr�R�W�P}򒿠*6Y���2�S�@,1��a��_b�6����<�`J���v0� �KZ8�p�x����"�Y�g��
�@�'�0j�mr�n��iɒچ����Pլ
�z�.��,]σ��a0-�1-�t��s����E�5P�>0�>�FRE������	Tl�ҝW������i32}�a@wy@�u��X�����18�ښ�O���^V�`>����BI�:B�� ���b����c}��<�v)��� N��$����z�	�,7��\�C��ZFVC~�z|�F��Zw$��s� �)�7���!��5�o�*Xt�1���-A ����LvvG�un;Q}	N��S���eRB��Nc�5i�C�c�;F���꘠7�a�������c�z�!0�}vTv }i��z�F��)�w�}6�m���ë�N/�ʢ7o���߰,m��U���I�ux�=�c�[���7���=�st,�-A�������}���K��0�� '����xQ���t�¢Cݢ ���#t:�/E�8�N����̦e�|ϱ�1�|4(Vhѫ<��<�wv%M	�7�+��Bg�s(�-Z�5��\���ʹ�֤�z]�Cp�(���7��|��n/}fi���Z/&Kg.o�ς9���^�Z�qhd޹n�K�ՠD�e��]��<2E��D�W�8�S`�<=���S�����4ld��Uj����v�er
�lH���r�·Ӕ���Vc>T�%�H�׹F�����0 ���u�?�.S�V��y�� ��z�N����#�ο(1�^-&���ݨ�����[�ޟ��.�S?�/j����aZ���I�c��-y�T���k�9�5�[jy�
V�t�Q��d+�F�%��@Ϩ:;�6|i���yN��)��ah@2V�oU3��)#$�BgE���t�<�Ѻ�f��;N��W]r���A�w�I�[���?�"I�^uw�S�Z��"�"{Ie��'Hd�'JC>5w�~j���8Aʾ���WV��N�T�X������Ia�=���%+��K;���|r�R�}�C�@���C�7�����*z���"�K֙�3�GR�����,�ȣHs����G��H�����*m�c|��zt�]Y�޹�n��:���%|��0�E�bN#���	����{��&ϯމa��e®���HK�rCgB�M��단n���[��S�;�rhZ�q�k2$�&�����e~1#����ǽ��_v���f;�����F��ݲO�e�J���o��c B9���� P����≹j�NɏZUIrPV�뒰)(�(}n�����a#� �e:4U�(�3�eV}�2AŻ��E"Hl��zsP����}��<�0�J�s��z;��ؤX���b�� ��D[���LiV���HP�s�:���E���?�۲������h��N�!$���^	 kY�nfA��NM��Y@QRDL�U회�{)�_C�H�wA����h0�(����rݸ�|"�_My�>������.�V�5��'� -����~O��o^��_�vX����Vl��;�jo����Ds���F�����'"Et�)�!���!��C�ܥ��I�p%�7�Oo��ŉ��y��
���K����W�>esF�fO�(l�����*���F-���'9& �=.9�C��$͐dR*n��@���Le2:��.Z�J�����$�ݓ�ɇ2��Ʋ�V��"\�}Fd+G-�7iTA>e�{a���}��9*S³s�cXX�^q�[���(��0�5e��ϭ r�馱�g�_ݏ�.�N�'B�G\o��<��L	6{!����_$�`���}��S��C�}`4�3���f_�D��@�'��W#��'��r)�E��2P��a�0NF '�-��?
��u��@kY�фD<��e|V7r!@tŞ>Y�V���I4M7�5��=u�Vi� �e�D�7�_�5�p�&S�(�n�Kg�4Ԫ����-���}�̩m�2刵����.7��65���l��� �K��i�� �5����uÐ���-��/���_��n�2�t���Н$<|QTu�4���WK���Q����˸���:�k�}eO�e4����(��u\)�Z������-��!�D�`�_	�R|��9�q�H��Z���Q�{)~�iw���Ǵ\�W�
�`���#b��Ɲ��̰���y΃8[m��S03pGLn��N�H,%��1��*]t�A|�3���^�Q7%�eMH�� *�\��u���C��M�w&�!O��~�zi��?���c���Oi���$�����N=�����J�JQi�1�+��:#�x<Up-���97���^ا���,�5yu���	�i���Ց�C.����*g�����"D�Z��:��"{�wk��$G��J�$�Ӵ��7�R�Ĉ�k�@8�i9bJVFf��,�e�xc��2�s��� ����iee�3 \2b�{
G�S������v�����t�V����Џ��?�I�����[k�v�Տd<��j.g#�����q����J)b�u�lLg�_e���.&�d���O%�J,��8���-l�]��7�����ݬ�5��U8[͈�$�Vb�ʍ��oi�0FvW�+�p�g��kĮ�KS�:��2E�rB
�
�,�@����?;�;Կ̥E�f�,�kY��c���@�t��e�s1@��x1���ʲ�.X�<sOK�h��%v���CyJe�8�����锲�/V�g�/Į�k��/�do����Bq�N&ۉx3�(�S�;+j��G"ҁþ��n���m���^�&utXn�K��aFv�w��{��>_�ۇ疟EPj[��_���@��\<6�"�:M�VӍ�V��?# �n�e:���x���
5���6��]!�a��Q����@��5,y.O��QII�8OZ��`.���������m�`��1[�7��U�����.{N��v���ms�.��!xh�;�\�Ym�a���1��/�l�G�j5�8�[l�2?A/+4ԤS���Z! �������&a����u���_p���D�(:�S,1�z&,do��ﰧ����'G���2UK�@�>��$����T��8*�)aGr�X�.޼,��B��o�*�߫]#Mo����-�A�fZ�aB�Pv����R`��K`�3
0hr�{��+�{D~(Q�
�(�䟖�l���b���%h샹ِ�Z��~V�Υ�C9���E!$����>4<?U� _a�W�Ƣ�x�7��e�}(e߉������h���.%��h�?\��0�#�0r�YY� �羺����}�o������:��*��U��y������0�3\�,��7oer��"�>p�9}Ĩ�b5����y��gW��u#ڝ�j����>��41�6t����9�kd_������j[� ���e&��j�kC��5� 팂ֈh�,\���9~@.��6Y|�0� �0J~�&!�aU&��Θ2�58ۓ;;2��/�s|jtK����/~z�m3Mm��}\蛽���!��]CL%�Kiu�uLrށ^p���eߖ���&S���ʜ�ف�@xBm��1����e�%]� ��TL+n�d������x�l�omr-��ٙ�Qnf�a�k��x�cu�R��鸋Rɛh�!ԃ8Y�,����7'�`���Y=�ψ��wH�7#�$��!��!�Ԟ����X�T�ͷ�y<X�gE�̓�u�X�k��N`���P�e�$����u��#�6�>�ӊ�佐>`X���@���\���n�fm4�!��msPk������¬��q���4��/XH�����ܟ"��2Q�Y����������$�i�;��8�D��V��J�K��9�< -5J���݂j��/Oh$�C�*��e��ğ��Hܫ?�O����i0H<%��qa�s��b�&�ӣ�|(��0�B3�:z������ Hs��Q�7i&GBrTt����m�mר��t�&!���c�s�i��.���:=�dD���D�:ԅ��s-�'��I3Ew�5�R*�͹��+�,�nV�X?�3*�NL�.(��&��Z
ܔ��K�$B�&o�,���!А��4: �����V�����u�R����k�p��[�Дj��������+qP��cȠ��k.?<�2'T�}����M�c��6�sV�n�z u�,�W���خ�����r� ��"��b\Fk`�1c��tk���l��
��=�t1QJ��ys�g��8�Ko1�Md�S�j*@�K#�!x��D�>���.�
l��%0[i����d�׬p�����>:�fT1�O� ��Ф�q�9d�.��r��T��ZUR�kȊ�U�z�e��ܩ�)�
q �����nGaS�J�*=��˱�=)�hً�w���q�}Z�z�.���|!1�����^v&�o�yG���eѨdӓX\�$\tg�o���ac��v�x4�K�����M�<�
�cQ��D%�G�1���"آ2J�� B|��E�X>�'���|��w��	�Z=�ؖ���%�v*�6��:\�OC�����ދ���S�G�L8��N4�Y�D��#���}�:g���0+�i�-xnՊ��X�
�����Mj���أx]�|����E���~pM�ԊrH��7w&����逄ǤGΝ�� T3��E��y���2�{�z:���Q�	+���
S�J	�GU�ٕg���i�c�}��%uo���N��Ex��4��3#�!,ɂ"��7��\!%����P����6�YZa�r�cԞ��ŧǃN�p�=�*EU������-�gF;�+0l�KcU�;Us�i�`"�#�q$�囫Im@��j�(ۄB�Z�.������%��b�Tq�m���BP��!Һ�I=Wҡ""��T��vI@6��9[/�zM��=��}s��y2�j�Vkf���/Lo��u0�>��h��E� ��������TF�t�ߙ�@��!�E��yg�3�-�m�lQ����e��ON��5E����\���o�[+R�tΉ�P�K�,������U
p���򑯏�0A���/�	�2��ɘ�>t��v[��4?�5����»��$��HՖ��c�\�3����u3g��f��E��#�*�w;p/� E�1�(�3Һ�����3t�H71n�A6������\�z�D���kU{�QV��xps~�E�8#���7V�G��:ZZ}����P8>^�c�/k�=�Ԇc@#2��{�ף��љ|�eSK��:`���냹�V���ʥRl@���b\#�/��˔�48�r�F�*e'�����֮f�ئ��Mn7��O�q�~�5�e�,���!J�Z����.eK�Fi��B�qO����LY#?6�_��v�� �����!�~D�QL�Su��3_������nPѯ,c+	˝�vi��
K����b��2Dr% lJ-J�o���n�n��Fé,n4&�c�=m�P�{h�[��X#�Ĩ�ёp���W�Һ'B������k2s^X�N�Q�i�C�Jn#����!lDY&���P��(�qY��N��!Ac�`�PZ���R�0����p�{�`.G�9���!��W���;��VQ���>�؂Jf�Ϝ�c<T���ƀl�DL���_J|��ftM.(��W����������������;����
"�_�/�4�2��A��:�܆���gDc>�M��L0�HE�t�r!VF�»�]� �KX�uh�JL:[�{z�p�ˑK�P�372�����9�wp��u�R����$��L����ӋɓK�߀Y�OJX����3rA�xk����<���+��l�_P�J ����*�>)��=��t�$�	6�Ӂz�w��8�mu���Q��Ԏ��}���U�T�D/�D�dŚ�彚0��J)s�J�^t��7�b:f���p�c�,����Lq����ٷϕ���k��F3N�׻>��k�b�^B���=J).�)��g�gv:gVY{�yDP�XZ���Abd�݅���F������/7:W�5}{�,���>̧����9�q$��ū!y�-h~*8��>s���9�1�������`ť���M��=���sr):yi�6�yBMl�=զ������r���L�>�εڣ��顶�&� }B�Ls����6f��b^𙟜�J,m4!�KL� ��r���o���o�lx�HIY��$R�C��W,�	�)��}�ż��͝H�����w
'��"&��b��N�97���3)x�d �v�_����.B���i�w��;�O�����?2W����x�k�?,bj�@:0���6��p���~YZ>��Cg�q|\���
nn����m���R+�Z���L�=�_
|�B2t�Q���&U*6!;�d(�i硇ׄ)F�'`�}2�a)�2�S��������#~�s*�ރ!��I���w�dX�~X�^��i���[���s���=x���=��w�,m�W�᠖H8�����`HK۳����gD�����1�ļ�g�p3��ީ?�?I��>�7K�lp�$��?�^0����*���2%�Lk3]y��`O�� ��oj���&��2s{:B~�;�r}�b�+n�mԷ0sJG�C��b�q������.�bH͇G�iD��v߶�J[��װ/	�2@���Fj�p��+��k��3���n���
�`��w\5��^4H�
����uPi
]�+%�h�K	�t@�B4�����t�`���QT1"i8��OPh�#�}h<���44I���G�Һ����ݲ3�ؘ'�xm
�����5�̂Bw����5��-�6Z��*��{���x	��-1�+��7K(�ێ�jKg/z1���*����0!ᅨ��٣�	�6il��֮(~��SV�8�'�&�4f;Z#=E���;�{Q�(�o�ҳ�iL<��Tｅ�nR_�c�����1=q�P���$]�,��f̢vB�d ef
K���(B�e��x��Hc�/��PS�Ko��k[y�N�qJ�5�E�RV�⁬���yVʺ�nj22b������4��>�!��7"����� �0gZ��OJ�0�(��c�q��c�f݈`H�S���/C*D���/	K�GH���O1���r�1�Ω~�g�b\��ӱU]wVŔ@���)ni�B]-�)~1�F=���/���=�m�?@Zjm8t�����E�b53Au�W��M�s����R)Éq���H�4v��ԡ�I�k�j�~��҃.�xĢ�j��_�U�l��,���&���Z�Ia'������lFZ��ݨx%l&�4H�b���'��u��h����ro�0<�.�4�)](A�M��2��m`�o� `�:"��e��=��m�ؽ�.���D L7�g�>a;A=�/K�i޿�l~bg��vX_f��a �^A��G��c&�R�y|����G�#��d�Ҧ�	��n��@ؔ*̚�̢�<5Á�fP/�QcG�&F~���I�1�m�������g�Yn�m/��v6��`��v�?j�f����i����8eS`��k��F�3���zj��kl���H��H��:�NL���yg��́�3�ઉ�Wj�q��7��B5
����I[�?���p4gޥ�Ջ:1��I,|w:	�Öf�j�k*#�HEga�js����s�w�������G(sZZj��6�ְx�s>��F'J0֐�M�R�������HM�O�H����>+2�D*�=��g�u7�Y�/��h�bRBo�yL	O��.�A�\1���z�І�fz�y��z�| K�a���$�){P���Z'����]��5Hn��$Z���.v�WЏ�qR:!	�J`�d,��2��l|�a�F���t�����x�8�c##xK���{�e�?b��d����PT[
.�B���|��%��h<�S2�"��˭a]�(H�?Ȧ2�ڵ�[����ļĮ�hJ`�q��K��/a��ht���uNH2�(f����E���|���4�Ӊ]l�/#䦁���Tc�͍B|u!>z����:���$�+�����|��ڮ/>1^0f���%�X�ռ�Ƈ��v1���	@O��T�)�؝�yEfD���g�p��B�R!�[/��m�:�{�?d�y[vf�B��ru�j���HZ�Lȶ���D�Up9�qv^�c�-��wX"H�܄}�Fz䒭��;�e\FB�A��L6fr!#�]u���qF�[��;V�BEx��y��*c���~�aZG[o��6�Bf�[�@�o�E=:t��#AA+��k��YP�n.\\��?��UN,B�� TR��fJ����8�4�[{>��c����)�(�&-��2�"ˤN/��M.�L�A�MS�e�%�IQ����CH}"�;��U~�oy������Q�{C�����������	�m��w�Nf�c��nN	7�3s��-hC�o��ªք+5M8l"���*����<�c͞#���a��p�-�* ��[��Z��1,z��e3'Y��S�F�`~��u�7�P�aFAAx{G��sK���SG|�����)���0�`a���l|+U����QK � �*Vm<D8-��f(N����Zs�JBc��N̈o8H��&�ۺ� �T�����!<0����!/h�GD�c��Qj��;+��S��d����Q��)6 ����Bk4S�N����X�F��@���ݹB�Mk ۹i�=T�Pw�qt2�q(���x�W�b��3�(y�0_��<w5ڰ�~"��C���T4�}����3}�ꪚ*(Z:���?��Y�ܠ��2�,<�]�~xݺ�����Rx���� 0�O+�,}�D�.��<<�t�� =E�����En����&��M�q�@�P7��C� �;�.(�ɼK,���@�*԰S�iWI����7�vr��w��o�SFj�Ia�U�Vڢ�'��j%�7E^�����r_N��I��OB�_H����a������Y�e{���B~͈t��T��W�h�Tqq��¤�i�h�K �Nhx�'�_���i�n�|&���{8j��͕���(g�&H��Yj^[Ǒ��x~:W�x��U�k�X�̈l�ؽ�ȳy�?)�����Տ(��bP��T!b�B@����O���*���=��C�7 ߞ��dZU��`J��Iې��1r�nD/K�Q�I�뚏2>�ss\�~2.&"P)�7H�6fɒj�;�`����h���j-ё�j������=+A��W���8�ub��8<HO.l~%�
!Ќ�^�Ӣڧ���6��%��ybA�&Vr�´�	�������7�O(�`�o!1���;�F��z��9�\p	j� �o�F����#Gn�����[��PD�V��0�*.��S��k�xAb�(�l�ښ3��L�>�*�wX��F����@D��c�/ j,��w�.BT=�D�ؤS�y���L1�|%=A(�>�r'A=r�A�Ս�?�?<Y�|�\����l�Q��
*>�W�v�K�L��)��sMjK�Z߁�4��\�\����c��Jġ������Έ㴱�Q*4�����[�R�sk���s� �N�S��~�5��H��E�hEf�����j��]D�Q��*'�g��Cb*L^l,���*貎�`4�*qXp��Ś���=~=���=*��&U�.I���x���%I���܃9�^�Ĉ�s���b3��k�B�����/]t�Mʚ����bʸ#�?d�ڹ�8w1���/e�Ȟ��s.�Q��� �g���	�S�J�ĵ1��5�P�[N�^5�6�����<���~n�C~�+	��4��qC��H�["�9=��A0raq�KrK�9�K�x��>���u�>�q��܂0R�w.�D��\�4«�՚(g��o������~��t>zt<FsqX�E� ��!`�&f�����8=Y���-�3������A��d� |ĸ�VmV#�v�w�2Pf੏�����R0{U������u�{0|8my��_خ�'ܢ��S��e��}Ω�9,jnV�x=�'��o�ԲE���@�)�2@[����,s�>����%�L�]�v��b��͓yyd������u%t(}SD���T�'���ڠ�|@���;��A��'�?>��w��zn�q3���tu8Ӑ�HF�hpAB*}����$�n�
NXG��������7K����a���10�@D2�)_!�Nם"�����Mk�A���� ��~��J�LeT�z�@PK�e�Q��+줭TP�ez��ص�K|�R�Z�
6xCF�B���YbxWU����1��4 �W���5�@�<7 <��A�� h���0S�()�0m���a�?���:Q'��-{͙���OXq�G�6����%Z�t�-����3[������O[�Un�����z�h[;X�#Fz�~��)_��qN�J�&	���d��|����'Itn���6{,AH��))
?�\I#O�y�r���8g�d8nAjл`VІ��:�]�w�{U�i(�S�X�wɥfT�9�&���*E�&�z&��Psk!�X}��	�?< g���
2�	> ݒ������ë�A�`�	?���=Srhù���`��RѰUz �5ѣ(�Je,��1s��2vǎ<
f�*�5N�Hq�t��kNLxl���Y�~��'z�V���@BB��j��$��ٝ�$(8�����kD;U9|l���g"��NӊR?�`9le8䈌�dĀ;#SLF��шihx�8�|�VI ����N�6��R̒x��j`>�S]�}���V�?iF�@���+QM���O�rt$@����P�m܀����A0B~
h��~7����.	��,�a���.���~.0C�q_�y{��:%:��FT k�* O�=���6�����,���)!�؆ܻ]JA�Ŵ%x�nK��h��'S�� y"���� ��X:�b\��?L��hF��>u�t��sQ�?S`�7��,Kf5y���A�$�NR$��@ӯ�b���r���u�q�[1@_��s� ,� �*�4-o� %��F9���β�]d뛸メ��J�cw��f�(��4^�4	5���Ȭ��m��YQ�؏�}��qh���JP�x�g��g �woT8:�zM�s�*k�(��E�Y3c-���Ӈ�-R�$6k9|V)��'�Һ�� �^�T8O[�{���+u8���C���Aw��ښQh�ğ���O8�*����<v�5Z]�I���e��K����L��:|�{:0�/��NU#��D��7��L���� �S������N��m��.>j���</5�*d~1�������+��Ka����m`�Ĉ��|Ŭ[��
ڵ�0�ɫ,���-���r'>[߆`.�wKbler�by��#�	��gOko�~�n�aT����a����I9��!H@c�Wh|�aOd�F�4�=W�w��(�I#.�w��:֝��v���v��N�G�y�,�U�nQ�2qJ��g� 1�v�a= �dD��� ��DL�*����pxz��������~�H`���b�m xH���CH%���i�.�[jV9,��+�2@D�$���jU�hq7J�CR�� g�=����$~�RLSA�5��~�L�mS�?�ny�<��6:�z3j�����Y�"�W�,ϗ���$��N`w�9?�J�I*Y���ki?�ܲy��/=�� �'�����[|���b7-�F�ߞ9��o�}vz��
���&�0��o�=X��4����?�3/^��C�־�3�¹��,��dk�ڮF��>�J�L�*~���������W�#��G)���ݾ�X�-R�\��Pt8��
�ԛ816.���>l݃��m���*���S��BB=T����n�u������i�݊�"��M�Y:��Vr	(��s�G�=�,Hú������9�Ȩ�g�;8JE�wǟ'i+IN<w��j* �e��x�\�K~A�����Q=�6�7_&F<߷���b��۹��B�b�Cx붶��z�A�?��0�0y�.�����l/Ua,�j:���z��-������Y�;޷������v����Z�8}]>��h�`Zmf3����`��vK]bMR���� ^�/W'���G:�$&w�ҳ�D��\�@p;���ckB&���E ���X�Oo�B����4��P5�T�b/��֕�2	�CQ���Q2��RB��;�Sc����������Զ���{7��*�!�j
<:ch���V$�t�c���Wxh힩b�n"�U+��`�Z�79���}��6������������/�0Bgx��f���e�:߷�|�Vk^�,�rU; �#��̻-0߬!�m���e�Ĳ>6���o��d5bd�6�_떑>�mr=�ᬫ�d�������%7�C%;� ur^�=�Ok���ko;+<�D���΂�����C]�$����t�^�]�3M���3'��,����{�[~�Z]�>e,�Qb�s e��,Yk# �)��{t7�m��1$�aT��ȗ�?���~�[9:�S�����!S��!�*��F[ّ7x���T[�t��_j�;;qx��,N��kЅ�E34E*�\��iU��E+3�UVB;%������S����i�L6��u'v�^Y�*� �b���ˁ���g�ڦ�)��ʱ��<���d����3�ƨj�Y�`c א�z�.)g ��>1"Q~=�L�C=9�Q+c��Dn�hC&n�IW�E��|��+��^=k������^�D�����G�c��ݤ�k,��%q�w��˛��3Ӛ(w�3����w~��a����ꄲ���T�t�:s>�ip���c��
�����~!��
����C*�2�.P;�\�<��d	
�6r�[H�8�4y��ۀ`B$gO:�0�Ӛ�$yM�y�	u]%VvF���׻���>~�̋�@�C��O����˲�f������v�.��{$no�7��B<��)n�Զ�f�Z��6b|C-/�4^�������f�Jbŵ[�Yi�d���v�	>���>9'�J�^0|g��C�  tLY��<'p\И��(�mk0]9�8i�zP:[Wm��7�ŀ��uA����4�0Xv�xʣ���� �*� W�߁r*U dx���*h�~K��gM|��ζ��"b#)o���rʡ��B�Tw�����)�B��,�)�p~��i��Աpx��F�qBP+���y ��G�������u�t�,��2f�%)v�H��];�X���r�_fo�շ��8l�p��h�@�>C�G�H�=5[]A�� �+Pb���_6�B��7?�#*I�V�#�l�/j�DG�Ѷ٠Oe��>�/mz�(�O�_�_g�AI\��ZJTZ�r�W^���9�V��XJ�0�b"Rbӌ��BܥK�uΧ���TȹkۅS��(�З�7�@W�rriyE� +��Bmɣ�B��umvVu����Ugq�[�c�ٛ�:�G^C��K�W�Ï��ϓ4��J�ؑ0�(��Uʡ�f���^5�4_�H^}����o'KĶ᫣+D�d#Y�+}Zú]�@>P�w�a�vv����ݎ�G�~���9���8��aG����³<�#��s ���`h��0��KFc3����w�xK���:#�s�Ϥ�$���d�|Z4��&�	�3�>H8j�bZ�L�5��&���$�r��F�}I�"j�A��TP W^�j��@ �1i�R�>k�4%1��r�]�{��j�2��_�Fn�V�S?]@�� �\�]|������� H�0���I�F��U���k7T�tAk@�l[���k��S�ԇ��bR8��H�1{�a'|
��wѐ����)�|�_�����nV��<]�v���Β�G߾/���Ka���z��A���"�pz ��@ָ�(�L#�ag�Ç�R���.�n�<T.>�f���व�7��»����ǃ���S�N������3�W#�"�;�Ȓ��DN|�\�`Lg���g͙�Wr������&����|V�/3�;�[A�8k~�&Qx����'��:$ˆb���h&Fǻ�,�OK�.v2���M��#I{X5ǜ"�?�qdh׏^Ƌ��A�п2/9��ܲ�Ba�fO�Qla?9}�5��}��]U��?Z�MX�j8whba���R,�1%�`p������|2� �(��b����!�r�ށ<�5��]m�1a��\�_�qU�*�a�JX~�̠` �D��a;\Lt[��dj6�ލ��߯�|��*����Ͷ�&˧�D�� �vɺ6��&����./�d���]�D�>&%'����-�׽~�V�j��ɂ�(�D���2���69z5�_~����v��#�F�Ӫ1%��N�cPysj��z�iz������p����� �3ڮ���%���<���;�Z�G�m�.������)Tnw�<8
=�	Q�������˻P���Kx86ܓLE�Pz	��`t�Ĺ,w0��m�o������{�W�>
ۿ���bh�xx��?��kӁ�J+��W���;�����MU=����M�#��/�*��_��~p}�猩[�#fvԔ'Q�{)B_
�l���[�^̭���$�E����T���!в�M��I��������a�=�sG�^3��Hu���t��̻�.����$��l�%��:���|VU`�*�z<,-ơF�ز�E��N{>�K�@�����눗��v���&�)����m�v�_ڦ��xlR_��</��������s��/�h����NY>�9��KI�$��ɵ�EC�[��8��U����-��;���d"��s&�寣�P�ez�$���t��&�a�ǟ[1N�d3�aςц�I$)f�Q4�\���%?V���|p�X���cP�&l)����x�e�C�zJr�7���H]��_VZ�N�uwL_����j���]�^OK{�����U5a�أ����"u������y��ap��=ݧ9Y4�G@]�CGl�?ފ42w����9���c���)~&�L�87�r��b�jS�Pb��7���lD��f��X�'���@K��  �qr�z��Wi�������{_�a�	�77^~��7_�ݻH���u5�?�����H50�G�y��ӿ���w�F���B����j����-RK~-��_(3M�}.����%#��k���U~�C��H�������vsd� �s���@>�����,���ʑݚ�x�`X������DW�Ik�:�l���4�LCl�����(ͳS�Q�R�Ï6�pz�pONl�4�w�w��BW���!$�w�7�Hfla>��*��������H���Tg�3x �����;~6((�T�AJrq�4{�E�	$��
�JJ1}�lQ����4A��� `#�������Y���<\hK�������뢺�g�\�Th��P40r�m��z�����=]6`�o0�{Y�
��0��� �������z%�?�wS�������nD�)��2���cO5��M�h�o��p��!�#�n��+];�Qǭ�{P��ʽ�����+���q^p�ZR����)d��=���"�Z�� ���L��/9p,-�?++v]p�����G �Ih[��Q�>�9�bk��pX������R>����x��K�0�Ɉ�d�О�H8�ĝ�ڲ#�]P�֨A�R�`�e���D���J�ڶ�ʲ�v��-d�|B��CU��r��3}<���I~~٫�]�tƤȰ8��`y���tU�T�"}q��>fU.:\+KK�a�b1�z⽞f8"��L���aX!%�+��8�o�������>쨋Ҭ�v�C9�����wN�0�0,e��L��+��8�5�X?ƀC+���}��qV��������>j{}?4!*!�>=�UG�<��*�d���ܠ#L6��t1K�G�m�� ��3B��g�<��"�$��}UF5Ƽ���������)O���m>���(+7�)QQ	d�7��$��T:�ބ��X���g�X*H�6�vBAL�w�ؤ	ǧ���^}X�A���3�O�,�<E��:�l��F�9�M���~�Hz,���T	 ��IA:�	�����y���rg���V�E�׹��:�ݧ�*�ld}�2�0s�Q��tg��!=}8�(	��Rk�M�~$p�{*�]P2$qD�Ċ^Gl�6$���J���Ҏ��+��d��6�+��RR
��k����4�^�c��K�e�\@���2�5uS�R��x��}���&~]��#�q� �˫��0CO�Ϥ�5���S���c���Œ8���I��A��mn�K�02��Hz����-l�6Oߦ�1(�����k�6	��} ,;�K�v��Y��2�݃���^sCt�:��X�ռV��'YٖFSp���@bpuN��H�V���`���׷Rũq�>����?Ok2޴����iLG,��L��֋{���o�-¤).(�e%����~N��g����Ry�R^��QXQs�i,.��І&�B���'`egw:�o#')
�
�/F�+�>��y@�A���s{����6�`.ms��o���,��{ )�Q}�fy�g���be���}D/�W�WG�d�-u4�e��#�Is���Ϟ�݆�k�km��ێI�Ap�y�w�
��S��(h1ca�B��;8�u�b19o�d����e{��?� ��k�U�蒎�qA��q��:��!g8���4�H];�������N���ׄ�5(O�ƨ,p&I��&�	����P���DAl�|d˚�>``I�$e�!�.0{_>�$�zs��Z|�o/��h.�`���n��+���J�����Sg
����ɉ�^i�
T��m�b�⡤SE;��R�^�yUf��vi��Ǔ�D�T�4������䊔e����$^��N1c.D.K�t��&%���e�XM�tՍe:Ŝ9-�Qw���߬vQ�l�a9���� n��Ja�E>�t�/�?�ꪺ��7�3V��A�?��8�q�<��/S��6�לJ| ���Z�8�Н��A|��o�_t���6�`�OG�v��	����͓|F =k\��|Y�>BX"�?=9�f,i��6���1�Uc��_+;?�2���S���!S�Q�X,����8�?�ߚ���;�n�R���`	a.�����#��A���OAh�.�j����:��u�+��Vt8�:��u���	}��6*UzDTҽ�u�ҭ]�*#�DY�y%���w{�p�~���J�Zt��%6�D�M�^GGrI������WM;����O��˒�h?��-�[c��f�-�z�"y@'Yӄ�ȃ%�w1G�tA̽��2d� >�sP�Y'�U;�W�;]~�Y��A݁�����R�J{��rO�S��wڽn�h�&s⽛*����8�Q��r�j	Cr��JVs�%��h���a����d��@@L��r	_� �:S���]y`[����g���-Q	B[&��ȼ�Lُ���ѫ�c� �8��>0M�hQ}jx[�C���d�<��ђyݛ*j�u��S*
��	)�ɻ�%��A8z4��e�M���p�s)A<,��y!2쵦�fv��ސ��� 8�Pkb��w5O�S�,[���يuF�>�>Ϣs$)-:�܈-�<a%l�䒆�w�t2�<Yr�F��1c��%���3��-�Gm�o�T�$s�H��a�P�Ĕ���a%蕅�D�g.?�����L�f9k��i����UϜ�d�Ǵ�.��,@�:{ߠ��j��a~� 3	�S$��er��J�X.D)YW=��j�Ӭ��}� Ȱ�����20֏
�ې���p5�c���� ���J��sn
K H���$A�y��'�w����eR������ȃ"}�*a�X�i��$-@Lw��,ֵ��鰱a�~FRS�r�J�Bb淪y�9uU`?_�9FI���-v%�x�J.�H� �[M1��oIL�:t�;���5������I۬-a��s|�mR�3E�$S���PN�畟�m{�ݓ��6½�<���货�C�v�E�^.�i�v��K}hiJU�Z���)��&�P��!O(�X���"�R�cKp����0I��d˓I���Y�<��>��˄�eJoZ�w����גu��7@��۹i٥X�I��&L3�;~��5�/d[,T�,��y��/�ie�+�ȸ���LZjc,����WJ������g��ߥ���έ��#~[;���ͿDs�8q�����On�9���wHZ�S)VBLayB���/p�� �1�� )t>)s�����C��t���ϤLYY�5>�i`�<��6Up;���YCn�?��p�MR0��7�����f��L��1Xdt��E�����]]ٱȏ�{鸧>���W�d�{�O�u��J*���{
]��2�.P`��Q���7F��2�3�1ٽV�I���n����BS � �+|�nb��Jw�Gkg����')0�I�j$a��ofeϊ�(�d�����(ҵ��<�4�� *M�>A�}��!H�m�Bs��S~�d�J�Gx)��ߊoS�d��y!�2g��2�mz��VGQ�~VT�Wb3���.�^����kn�O�sD�[�W���y݊�I�U�9Dk{�I����H�:�CO��ø�h�����y�`h�U�.��yF���x�����,�PL�-W[��~]���
}�s&�x�Y�[�O���`!�b�X��/tW���C�R������P6��p��� �!�q�~�rWar}<M��u�v{��݇E�G�}-����"k	g�/���̹�	��>�T�1�{`�rיQ��ζk�����Z}����0H��̲d��c�C<C�|!�'�<&Ue���ǂ^�7?�NkO#(���k�=�=[X(u���ӝ
3a{�Zn�Ϻ`�;�M�����*\�So��P�"J��kKh�ꅕ��U�7��&��w�@�Y�_cs0+���R﨎&�f���{k���G�:��fT]u�Q�@��f�+F��[��e�o�#O�a�������
8 >�t��=J~��R�|}� G6�V� �N�޵K�r��	���X���=n�ea�����	��7?��p~�D�_nl���>#���%�S�Γ�u����.>p��������\C�4��^��?Nu|}��B4����W��Y���H��.���5G!]�k��`{�I����IW��_�h���N�eǅ��*�:����ɋDe�����?�2w�7�ք��<�����xc����6嚰I��� ��s��6�%�, �)�A+f�:��@E�?��6�Bs�Q/_|w����ɹE��Z�y��b��H�a��#K��08��Th�]a�i,f9��[�b�"��4aZ�8"�t�go=-��ͽꀐK+�υ�iJ��5�����\��nor!���'�<�ɰ��"�10��c����X����,x�K�w�U �4t&D�P�K'��V����DRJxz�'F��k5��}.�BZL4]���|z�`:v{��1g{9�/ͱ)�d��hI4�$��f%�M*�	������N�~.:�gp��S�S�Dj������N�^@d>�	]���$�H��)�,(!7�#��3�4�hl�H)�<����Zоd�ao��#ST�yȁ�"|BL�k^R���j(����rJ���b7�w{:��&�/��޽����8q�c7�jҴ������B����2�6�G��!�Z����>��XR�$��0޸�'h�Q|�I� �ڀ�Q��aei���4���v�&��j�t��u�nv�_Ϗ�˔�	F��ue�]N����m�E'���RB�7�
3��	�}����
����9�:�!n.Z�WGT^�w���!}��p��ݘM�l<�5M��4_x,ER���]��h�3Kz�#���Q��
�>��2�@]E�q�YoJ_,�%hq� A����+<�9�4��>��-��d�bB�v犩g�����rp+�	��\6�
��G�}�Chu�%��U"�e��|I�o��yz����R+[G0p�y^�������t�yU�h�������,��N�'���fQ�!f�G�N����3�6]�u��7��;�6��d���<�(�����y���V��I���{F�x\��K�͋�%������4	P�_����S{���~Q�,�b�ۧz�W�����:�>M<�������h��I��}>��R��`e��X�U�!�,��f�S@Bo��U�����{�S��l�X/�Lh�C8�j35+$�(o�IF��n~j�^�l����r0�-^����hޠ+��'}�-�]	ӿ�L�������aT��k��+�X��:�v�ed��,�f9ub@z��L�
iNt�|��Y��Q�=�a�7���bM��aei�ʉ0���]�Č6Z����	�W��Ķw�8�d*����$����;l� ��xe���?P]6q��9�4m9��)���a4�,湯�dSl=��&@�V��]��m=yx~Xt(3���>CZ}0��\.2{��2�ugj��x��N�VK��HSϞ���H:��n�J]䢌w�M�f�q���caH ���sooXjVWs���Z���}_�����xa���[���`���q2�P�n[��6ˢDu��� .іֈ���G��a�_��:C��Ud��k�
���`���F��R2��yF@X�z��h/��z�X�9}�����طT/ړxo��՘�IyoK�҈-(�����n��x����0�2���[�k�,��Z;#V��v��@'p�f��ZM?���x������?���#�+A��ߔ�N�t�z6�f�_C�/[1� �逜
�����58�<c�fՉع�i�f�I��W���L���5lZy��FAc���;t軶�`w�Z�`2e�����/��b8�3K�9��/}G��bO-�P�A�P�¥Ǆ��6��N;�^� [�6�M�)/e5�E����E[I��P5�����Y��	�x�(�F1�-5i�"��<��"�V<�� �A8���e���y?�E�%�o����k��r�D�j��C�]�dL��T�ma����r)ǯܷ�NO��r�CN����~C��R�ZN����M�c��20Hg����0��:A�SFIre��b%�!�f|mᶗL?���,�]Zֹ�\�P=�N�~�z'Z�<�AM���.�}���!$�Y�n��M��4^(�3v�����Z'I�+�d��4]���K�T�ğ��THOz�����9�r-z���e�C��J�~�!��9���M�&�ѓ��J��
�r��φ�|ù)/!�Ow���
z�9�e���`���+��7����k�G�{���v��B-��;�3�1X�����'��.䮫��+c]��Vb^�:��s6��	���&�w@;\_;1 �$a�KS���,����W�$�-��v�^G�f!t�P�r.z�y�} 
L�k[��7Ϭ���$PuQ���D�~�W��R�ṣ�������U�8[���1`q�x�]�u�@X�P�Do��*"UO�K�,�)د$��m]'"���ʇ���0�b'{����t�&���)�?�q1R�f���Y��� )���I=��^�f��l~ٿ/m���v>>���1��7�d:J���7e�g��[ug}Q����׀��fീ3�&�w�.��80L�CW�Q?�Ye���-�r��U���6.;��#��9M]-��X��I�MƳiwc�s�N�c:e����|��a�]��@�����=]����O��]+�U�K4������d���\}�`5��
r��m�{O��Q
�jV�'����.�{(q�T��7A�,(("�d
-y�˗�)1�V�C����w��^�덨I��G��CBb$%��M�0W�ѓ8L0�.vrP1C6d�溌)�� �rO)�s+�0��k<7R���$
p�Ε���j&4��������5eF�^J�ʗ�^e[�P-��l\3��<}b� ���E�$J` UMU�ҧ(����18;J���~����rE��2O�����yּ|^�AX�R5K�Yc�ġM�6&A	Yv��?{���$a��0d��ܞ 9�C!�]�us����:�*&����fE���1���8#)�HV
,e��V�;����%��q��Ց��SFf��u
=��v��K�ulO,�����Ct18!\��b�g�����*�6Y������(�M��-�dk��I� �vX@Z���|ByJħ�U%�gU#w<���X`��_��q�I��6`��bќp�+�������;�a��>�?��� ��]�d�����G�gS9v)��l��hqj�(�zN8��Q�[��DSٺ8�m�{ҍdg,�4��xCnǢ]:�UE1(��;��Y)����Tp�������]1�1z�}��BT�*��/}z���5�s JRh�E��uH��a�Y=]�qC�Hw����D7���{��/��ݏ�N��H�������lޛZ�:~&�Ï����a���dg��g�sfR��u2�U4�mũ�L����C޽�d��,�(����+�s8�p�`͖{���{����Ä��j;@k4��8�6,'*��О(p3ߥ�2�ֲ��%��Sg\�O܍}������G�[*y�d��y� �bk%ƶ����c8�_�+'	(�N{<�1�˰c
����!zbY��{��F�Z�Q�=������ =<�����r@x�':��V2��us�=V�u,�3	V\�$��Z.�̚W}��L<fg��뜤`������f�6Pa��#K������i����g��'3!l��Ё�P{[P��OFKo�-�ҷ�ú
���|�o�7��4Q,�}�g�^ �9l2�c��������T�&��lb�e����!�4X��:���a{�g���G�!{-Q���8���ch�^���Jm"�g���w�ٌ@Wt��0α�-q�PBůW�Bb�]���XԸ�R.�!�q�$����6gqq˽����TÂ�L{!��G_<�%Q�Q�k�^���L ���;��(Bt�#���&
����!+�� j�e�[{+|d����qN���i2��B:e� ��.Wz�3����L\�;�����bW�o6ǅ��b�Y{��-�	 "U�Q��it�)b�Oոv�c�;��ܔ>l�ݰ��Vٺ�&3T��R�Ũ�y�=H������,���z��"�*�U�������fbmꪅ�J�`�uB�+4�S`�P��]@Hx��Rq3������"��"0��������l$�%ݱ����.��~�~شZ���ӏ�$�{92HA��$�+?X�ֶ9Jٚ�d���kiuK���T��w9�&^	��˰�Ƒ���	󷝔��;X>OĤGGגR'�.MK^��ZQL.+�H����:�݋\��
Y���[
���)��>���:���>b�c�-'�ۈɥ��L����Mх���NnR�5I��b�>"������⭳^q�V�_���O+
�w��QwD1�4��bN��������%]�85ɚ�-,l���O�1��j��7�xM]�c	�k�
�|�Ս]˹l�Y��pY5���ey{������.����_܁���lL�*����	ĩX3p����O�I�gXgp��,�m��߆3��'��\e��H�_��|l��:�@�CD���H0a-Cu�wiO����|`}Đ����9�h��)pU@EN�v�'h��kCb��"�����ĸ����v�p!I�PZ��(�%�Cz+>"��~�-1��H[�jl�mk�14�k�1�i]gt`P��2Lx��N[_R��3Q�U��X�=,�jBF	���5�W,g���痢۳�ݵ�qG�QvЧ�t��-*.�G�~�X^�fꯩ>�U����T'L��[���/OS>�yo^,
�C	�rQ89�gd�/)"AA�'eKr}HU��a�&���E/����*
0a�?�8&]�2��G�G��7�=YU2�*�2�M�؄�A"G�j����k�D�")����Xֈ�� |������5�O��)?a�u�O�`�HD	5���$�1bǤؗ��D�="%�+ɸ��3	.-�S+N�}GX�-��Y��F�ٓ�H�l�PQZ�=�o?g�f�1�L����y%�˦M��;�c�*-�^�Q�M�{@���/��E�h�5Y�FjB$S��eHs3�G�.�[�d��/2U_�ܱ--y�������1l����[Ɠ��iVU<!͑��c;'p$7�Kѩ�,��;{/4�F�!Pq�;�������U<*1A��4�#�Ny��6�j�hgP����>W���ow�.a(Q��]E{an�KHG?,�7�R��S*#����6%[ˤ��������z9��AA�r�L	K�H���w�l'v���>f��)�,���d���5��v+����\z{K�
�X�J���3�KY5�M�ٕ��JٸkK�	)�P���@���鯿���wɏ�j�X<�G�x[�p����>?3)~h���]��1�L���w���8l�6xhx62��!��	:*�zW��	$��l\�(!S&�!n���������fJ.��o6��NE�D	c-��}�gRL�J��5�M�D9=�"TY�X�������k���0����e׽�`mY�(���sqDu���2����2��6'}��)��CH� v;��.f#q�r���ı`�(8��c�t~�£nP�ϓ]P��?
~��)��V���.
�܃v;IU#▐����A�Ӡ2�^�(�(m�X*�'X���Sv�D88 �X*�h��=G����_h^Cn(�H�a��C����S��*�<b��닉 �:ִZ��>�dX>��a����� _~}�����9����o��H5�1�q�IX�CK!n�%'5:l�s������RF1�ncݻt��II�'?9�n�3��#P7wLC�%�Vin�"Xu���*�bϠi��L�dLl�1/%�]MS��̺��278��r��ywz[�h��wv��I����1Q	���0>E'�K�|��_mމ���b�'�Aƽa��2�;e힭�����y(=k�&N�{��l���jqWPT*�Ơ�|�����Fz�-Ssb�IOBh���{��C�h��.�y@G�E���.}v8#N�ý���z�)�N1 c}�3�Gh�c�	�pq���[��.�4|�5�8��<�kZ�6�E�A�pw�n��׫aZ�ӗ�x�������/�c>XDd����[MS��u+Ôo!�l{�����<i�T�C0�<���}i760 ��&@qK��@�H1����h�f��?k��"������䍔,��	��\���L��G�ͮ<�h��<6�Cկ �C��c��T�� � l��b���i���5$z+?d32�G��5�N�^"���Z/�4���DL�G���n�P��K���
�?��}c��\��hG�z#��5�ҽ����,��5=*�2�*� &� y�S���N�M�kNeL(��q@�(Q0H�6t��>�A.�N�3r	2Q���U��b���b檱Ɓ�C�K'+�\��k �fsr�.���Ŧ�	���r�]�Fŋ�xb�X���wPJ;獄����k���uV��Ӧrta[,3Q~ʦA�1(3�jz+�:�1ye����[��˒���s��8����b"�����fԑ+��}�4���b��� HSs�#�n�P�p�h)��nC<-���F�O��$Z��'B�ז�da(�ܦ��I6��習���o�I���zz9f�����խ$y�@��X��~��T�����W��E�$��^E�v�J3�Gwy�3��"�H�{=���b�a}�J�Cs���������t�EP]�ko�2�����3�uhެ�c������߾f��?溊| ��$Owf����LN�Jk�ȏ�Z�C�:��adȏ��O�m�|D�Q-��w��nl ��Ƒ�f$r�T�h��K7"��,	w�@��d!��SY }��y�$r�:X~�.��� '.B���y<���\��УT�9��֯�o���W��&Se�r�����b�l^����V�~�^�X_xh.�#�Ǽn�^����Ԩ|�w��a,����X�����k[�;q��E��������P��3�%7�oO`u'����D]���dT�Ū�т-r��p\!jΏE�ێ��Ǝա4dZ��	*Y�3l�0��2�)�NOo�K-'H��4����:��UFQ,mu�S����.J�m$�th#]�.-��n\�d%��(�O��Q0d�?�C�,H��sf�>����K���F��x��焟y�tq��Q��=�Mg���S1���?��_f��~�"������0ҒF�;�ʥ��?^�lYA���L��`�m �/�U�� �OA��4E�}�p������]�C�p�۫��PT1S �vE�Kv��4+�n�[�1T������Q �;c��P���ud���������}�f�YK
���zf���-��n�sJ�c��.����w��I3e�ƞ�-w���2���|�p?�\�y��,#VT���	�·�vEԅ��@�3�A��Q5�jOT�L�maܖ�@Mp�\��-���5.$�j�C�h�B� ��ܾ���/Ǒm:���8�߉�m =-��v��:��1�=
�6?�Ż~��3E�ݷ��8��M��B���������G���#rǀˍ���jf�T_&bY�o�6�~�ĦA�hn
^R��r+�l���ܵ�^�;�L�G ѮW �8H��=O��K�[��:�~�z�L�4/%�$��ު[J�M&~��i��q���k�"��[I�9�" Q_��3�9Ey�D>L����D;����@^,xЭ��2���N���;���[�h��QumU[D]�Is��Ӧ	����N��_.�)��o:I&b�f�����$�(v<'�5�9�y�A=۽�w���`�������WLOKмrt"p�SJ릱���65V�$�����%�h��3O��/d~�ZT\e��eoDB����A�S[	|�΢s�s;�;!�(hD/~�$�A��?���^?JH���%GiW���[��pօ���C�Z�If������ʺ�1�%Ɇ�X=����f���'|#2x����W-�ʊr���"W2�6��z����#g���s1-�a���5A�9U�J�����{I�E=u��*�4::�lq��������Lh���c3c'����H�^�{V^���6[~v� ����OV���(I,4v�%���w���������.�N��+�U>@����4�]
��ȵ��#3�d���JWy�{�:� ����m�D���y�)�>^��|��=�3`P5� !�)J�'�� Řϵ_?�U��u�}o�fA`��£����H�������h�s��g֛t�R����V�n�a0?��vL�04�{E%6G��$�C�o����I�8Kv�c\���f�Y�)����dC�H��l�Z��Ǧ���}ۈ�iY��q�{�s޴*�^�2�
jd?�Y����L]�g�/4}˂�ތ�</0���q2�΍͡MF�������^�գe@9�����U�2�v	��C�\��f�
��g�ʫ�n��b�i<���}T�m�:N��A�DUzz�Ti��Nͩ�^윶��`�	l������Nue��T�sY��������y!rX��.D�km���=(wO�|K��w|ߥ�Hk*[��\�;T5��f ,�ل�ך+�!Du��?�����Xu��� � �IP�<���o
��8}�3�K����)d[�x���.�;(�� 9� 5�����<��-R�x͝���+r(��@�ؚ|5��u(�s1nN����~�-Uy"�z��e�e8u����6�sn#�΍�߇�e������t����4���Bx�\���$��&���*+Ƶd1K<ć˙���#�!7
,w�DXԵ���=�/_���K�e�%㏢]
�{.PA�K���H�u%\iOoy�⁫7"
��7\S�d�XE��O�\��p�u6n�0��%莯A���I#�Ϭq���j�O�E(N�G�u�s��R��L���d��?5���3Q����e;�����tƝ�/�k-.���Z}t����;/y��ƃ�ѰL�_$sJ���zb�k��!�h:�Z�k��X�y�߲#ij3��,h�_��*�����􎞱%<���W$�l�p\-�k�[���u�J}��p��f͖K[S��.h�B40.��Aѵ&!�h �2��CNy���iC�tU��zΖe�A4�ׄ�>q�������M��?)��E_xԩ�Pɪ�CY��W&��H�%M�_W" FGv�M��d���V�MiyyvᑚID�� ��u?��B0�Cy��T;��v�l?�`��J��?�C�����.߲̳���e�?�sE�0+]�)K�DL�^2��T��4/Ex��Y�1[��z��VW���1�})��_ԓ�5��@ȅ�8��3���_�&d�O���V�b[+�\�����#�ok�Ѻ&�-I*
��l�ť���5����T��.��e��J��KŇ��2�j�YD�u�ނ3����L#K�_�;j�ħb��|\N�V�.O�����9�Oָ�����l����rb���O�.S3./~�Q
}�9���HCawR�X���!���C���8�8�i�%�I���<�C�.�g�D����)�}�W���G���Kfs�$�=��`3yt����82Q��=d�ڌ�`՜-lqK}��b�SS�z$@��4���r�9-	<28��V���L��r��]z������<$��F»�f�Oxʹ�8�f啗&W#t-�0(#�SJ-���r;s6������\��Z���㒡@l��!������N�.���<�K�7�N-�C`���B_�8��~g�ӄ�0;+�yp�1\J܍A���ņ癨� ��@���4���:�|>���췚�����|Yi--��ƚ�� ,����uT��r7\���J���1ob�S%�E'Ҵ
ի�S���1��"�<;�]7�+RW9�}Y)L�B�  [X�J� ��1�Gpt=��Jj�G��JhI�B���	Rn���_u �Է��z��;��A�n��t����f=�~5;L�ؿ�Ȇ ��*`�B8��5�2�4 X8�<���P���P>3�.v�J����xr�Ҹ�/�� �RDMt�!�)IS�H�]�|%�*��pz{"�We�^�0�MEAB�O�v&��C�K�y��$$�k?����A�E��m*������>®�5�q칂G���.�	#���0��#�Q��d���ǸC�ղ�l>��ߍ�����VQ����C��O��� ��o�X�`P�Tj�}۪�4����鑍��e	�},���T־�ڄ��^����'�o�-���$��7����[�q�ક%��Y�I>*d̱�+�o(�\F��_�ʹ�FW�%/�d7|y���P�Q=C[t'��h�g%���?��g��!�I�T<�jz�Uc[f\\����vI�n�+#4��}k��֊��K-hp��
�E>�纹N���6<�qv���:�Jlڧ�Ĝtm�u�u� sx��UC�&�߆	>��&��#0Ghf2��Q-<}�S�_*�0۸)~�7kB�VP탠n�ۧ��/����-3��׸ROKQhH����y3�̈a����3 6�g�;�_br��?7�DS���A,Y=.�R�
Q�����Ir�D�ۂ���: )s�,��u�?�dw�$�Ta���$�R��=��ę���&� �)�����/4;���Yx�M���^�|c̶J[9 .[kw)�uf�`2PU�ҽ8P����HQ�ws'Қ|t��#/���p��U�M�u4/��d�t�����|\�0)AՅO�VRC �P�����aS%�d·A�7�e@V���&�Mp��M���bv�<]sM�+���F� Lx�{	/T�0������h�I2�Zٓ�F�Ǆ>��8�7�v��w�
!�oܹ?��򶚌=�_@���hv,Lo�%Xf�^uu �L�����&��Em��s��B[r�J:%�fÃ�.8V0O�^$�ݸc��)�e�@����i��9,��Z%���Ķ��!�z�o��I�i�JRS]�NQ?U|˸}���nh��6��6���$�e��b*���+����e`�F��U̶��V�ư5p{@Ȉ��Z�������gP_K�1!H��2�˽��x@��B���=�,W�=��\<�{�%B�@ �~�Ϻ/@�?\�nH+��!`\���8^���&�!��C���Z�d`F��cb�����������Xq�X��_��-RC}��n"'��bF�x4osi�>�z;:��Y>�%oK�x�ݺ#�_�g�M솚������#7�*�R*�z����
�i���^<t�"��oT��;>�vЪE����&~\𼁖�b�jH�oN�\r��C�'��x"��{�2@�1�����;c^ؓ���91�w�԰�y����ԣ`]3t��A~�r�S`h�1��K�?`;ӏ�ӬCgVd�_\��C���8*�����?)m3?�仉�ߺ%�wFjx.e!�.�Z�5�Ӛ�Ӎ�b���G>�z��8�/�C�GX������1"�uۗ�h���e��4}f]1���򽑭��ڴ�z��BMze*Ƙ^���{�4BX7c��!��עQ���c���z�:~Q���;,m!N6
���w
N�xG����&ʹ˗62aZ�l��2��"��Ij*����&.�M�?/��N��5'K�k�L��J��C|˕U�����^Zbe&�d�� Jvk4��$b6�R�#��C��@�d9,��,��֋�1��i=�V���6�r�9"���-�/R��G�2�:�/']ʨg�`�h�p�p��ϼЪ3��s-��[�K��xR��X������,V<�7k��ѭ<o��e�s�捷�wko������_OpV>�_��o�x�&FJl¥g�2�b
����9�����Wq&���t.1������b�4<H�j��e�;p~����_�wQJ���J�U�_;	[<D���E����c֦����Ą�˓]Z�p�W�W���{�O�3�0����J*.�!tEjn�_���2�O�̐�;�]ɮ91�/w�'��$�n4������\�c�c�1r�x��V�һ�q���Ptt�к2)|C��-KQu��XxtgB��{GN��ԼM|:G�ߴ�"��t!~݁�O�3[,�c���c_���ަ΍�Dy���~@&m���#��!#x��K��=�����?lt�V'1;�t��̣H ��(�(�-�2��I���#�Z��F7��ޔ��y7q� M�p��,L���u9c&HEԬ��qW�)~����I[���o�%����\����7�<M�)�W�a���~����3�1ҕ����GMKM5�c,{�r� 3+c,#���[&��"�:P��j���Q7�Ǽ�>�� j���V�n�i�A��s�V49�����.���:g,������u�S�� ��ۭST��������w�m�����j��f��,}��'$ ��U�2�~Y5n�Λ���ޅac�q��	�؈�3���r�0�a���+���UI[�'��b]�?�,�K�{ҏGC���{�d���'Q��g~�l��E�^kY9�/?����d�d{}�L�.�kJ��叁,l
��ҿ�7'n�`�{�_�\m�T���,����jʏ�4먰�g�3��&{}�b)��#Zʌ���.�������Zf�Zo�Ɛ�y��}�8��=����Ȥ6J���X���oSt+�\n�i���~C�0�B�ҹU������xI5�W�A/��o� �t�c����	�?�����?�x�ii���S��3.�8��F "�:��qSѼ�I���T|c���]�|�pHJe$7�)��>Z8<�?q^Aek��0��<�Y� ��X��mW�h]�@#]�<H����mk}UYQ�ѹP������?5j`�7%�Q��X��
�"��'������z�ܽ�<��(����w�
#J)Dv���*g�AY@��RE���H���^J������Er��Wx��v\3���pN]h��uWq�FgYF��.!�?�i5����"�I�N��J}0���KN8��ZkR߻����%ѫ�/KHݣ밻��t�w�5���Am�����	�f��Ki�8}�Jab6S��`ڟ!�s��:���*��;U�y���tJ�������r񬿠v�c��	��� �a�h������P������tv>���g�<:���K�INB,Yj3$Z١�-�f�u��
M�MB�e1��Vчr�"�ƨS;����Π_A9=����aΎ�f
���	�c�`z��p�d��3��2����oX�U	֒Y���S��SSF����Id���?�f��
/�2���z��YbJ�I�)�Ø��$̰JL���`Bf�ZƉmI��:���˯��]����_���B��D�aa?�A���k�Y��gE�� '若l�=��v�?ydġb�U|UU�9�݃u)(�2Ph1:��s�鞐ewm��rsO��!<��(�摳�5�+Q��^C�j0��O}�����[��U�����p���QW� ��Ty@:��B�����B�-@5N�wgd)����#��ݴ��[ՙqDOP܃�����^E����-ܡ����[R���Π)�5�&����ȩ�qs�%?��ܦt��Zy����
@�����t�<�� �7[ha�T!62�����
�>c�B)��@��X~��	��Ck�D	���j�]Q�)1v`���i�,��A��I�#��Z6��o�1�E��/9>�4�����twqnY&r��/�c)��v�HB��y-�g��htyIsYG'K�XR�#��Iߏr=�:��}��1��˦���{|q�����DI�>Ow��bK7`������[��g9�@��&����E�f6j�o;�n*Me�'���j}��4�T�j�?�k��V��u(��K����r�۾H��:�~�H)J4'D��7�{8�`!����{~Ȑ��I�Fh��Ĥ�:�����x�fyv�xN�f�Ԡ!���m�K�f��Vʆ����y<��?|y�gA
���|ɧxTr���a�{b+����~�I7(8���O��sĻ����Z��h�r�]^Z����P� �������1�'%�i�G����5[�X��d���G���
׭�g�� )���5^�������� <�4��E�2�+���1��ZZ|"�-vh��8��T�j�J�w��6���*M��a*�*��h��؟�������o3��X��:�*霏^z�=ά5]Tzfpz�5��5��k:�:�����0�@���^e#�U/5�@lx�9#�/
�)5��#aB2��|Z(����	^�!�K���v�d�U�7��BNs��Q�������K�����7C��pG�F���jIj�b�E=.c��B-5����G�.�%�:��9͖�&3|H|Y��� �KLʤ���<���9�gc'F�s�|V��Y��'%ƣ���{�@>9W��bQ�@��	�����B�7�9$���tOͽ�v�����1���<"B�X.�?���!�����a%�<��G3WDȗ��a���p��Y �������=G�y��`XEY5D��S��/��*#�2f��4p�*��c�
7�Ә2^"&�u���n��h�S;�O������t����"v�U�3f�I7/�/��^F\73��7rEaZ�6��׹x�;b��)��jN5�'�л��eJ)̸�y�C��s�*�x�_�u����%P���s��-�aMc"���l-+�}����uq�1�z�f��Dm|����2���?q���6�~�u�g�\��m��A0�
����i��˞��~�/��'ڏ�/� �}�G�e��d�ϴ@z�FMR�"dH�My<Ju��r�������Xp��9Wr5�1%29�1
�x��B%���tS�v�Z2d���Vpԍ�%̨�>h�G��I�#�Cs���[��L���k�K��� JnIo�"�A�0�G�E	�[�K܆2M���lo)��@W�c��Jf�@U�$	���䔋��۵�������OL��M�?�M$�|�)�f�x%�&EQ������>�\���|P�SyQ����3n]���rKt�6>��ѵ�j�A6��t5eHC��������q����=q��n;�2���MMnb��<�#�Y�n��ft�;ЍH.]/^�o���Jxͫ�X��|��i�H3��,.My(���S�c#NĻK�&���Ǥ9�s���Ӂ�8<=
0���m.xdr]lh��Λ�9��l�zB�^)�2���A���b+�:oѥob�	3�ȵ�)~M�F��"��$�VU|5�F5\i`0~R M+�W���sz�J�U�/9��Xep���#"�2!�,}ϣ�p���������b����X?�O�<O;L��&���:>�)?7袡 ���Y��@��k��A�X9y$w����d�V�@x�g���RKo<5��t08�jzb�%��4�GB�&�tP?��O����x��Qx���@I���=g����%$�0����yC���4߯�%	 Q,�ޑ�Rg��[�le~�zvM��~{Ce�� g�1@�g���K3��dS�+��m��^�Z�
1ދ툉5�U㸵�I�s�i�{l|����#���[l$��bإ�F��0Y(��L���P����E���&<�k�0X�����|��IoB.[��[cDЖ�s�/:G��>�sZ��<]�,�ºz�_s$7B�e�E&)��Dv������^�U��O�0
�f�[�t�k��� I���|�����'�H���l�0�N���_���XZИ�[�3 \�.�u��Sk�峨����ѽ��")�	�/�5�_p;o���ن��4+͠��
���5Ě�g�#w��C��]_*�ğ<e��g �Pw:�Ť&��x�'m�����O#ܘn疲z) �QP���>x�����T����*�IY�4�:���M��EOЃ��p���vPJ&���	�W��@��'
.�q�HU�{﷽���	a��u�M��S�d������Hk�eK���O�[Jb�QCc���U�tm7�l��Y���$��C�o-3Ӳ�B��`�q'Xp��oN���PA3�˶=��Y�|���=���r��F����m~�����I9n��6�.��B��fJ!] ��!�Gf��hL�ZǢ����i.4���@?z4h=�;O*
$ ���i�䪎ϙ5;��{)����vv+G�p]	՘g�
�u�3?&Ǡc��*Bv�B�Ӡ�0��.~+X��m���Q�m���ߎP�}���쫩��BeRd�F�B��$�@(=ܫf�����5G.��#z�0-n|�~C�d��ծ�`��Tv� ��8<�m��>����L��S�
��' 1��k ��_�M�m��K2�>6����< �D="��x�e��٬V��lS�)��2wZ���$e���_�|�	J\���l���k�[lB�uO�A��&�l��^lS����Q[g+�j-������II��",��ɑ!�� ���y�&7;�N��T��Կ�����>$cQ̐�wI����&R�V��N���/me�Q�Ζ����{n	�W�����<!��4������Sn`���C.$U��3�E��ᡋw#��j�@�$��e����z�Bj<�ށ5Cm�2�E�Ǜ�k�X�Z\%��������t�������0�j����~��1ڪ��kҥy:�����A~"�x�/�n�Tx�l�}���1�EoQ>!l�f���'�3��ǀ�{�(!4����c2yk�t!QKPc}�=?J�~�
���n��\��vM��̩��8�i��vb�^��>�z�b�S��K�}��.��<טB^j�������⨴쪑��hl��w�!:2���6��s~e�}M���b����Uݍ��|�B;)�ʧ��_��� ���H\A����H���<����:LWP�A����v-1��9n�D�ӎ,�e~�oÔ�a�<�r������oyQ�K��|���_�tJ�1���G�*`73�6Jp��|��6�n�2a�J�� с!�a��N
���Sd7{ˋ��l��(�EIp���Q:&�F]�Ǣ��U��ܬ_
�F���"Gh����^?fle��pkQF_�N�D��/I��'��@K�[-�&�|�����m�h)r�Um*:[�p�I ݅ܟ]A����U���b�ފX��_�;¤������l�VɜJ�k��[W�Fl��~;K�s1h��B^*�ȣѾ�ې��\���Wy�'Y�O	'c�VHB�	�)��%vb�F9���̙ۜ��$��iHH��{�/*���#��}K��0T[=���>��������wsO�yµD.&x#�'I��8���%��,�n�K"�p�[���`��=�]�8Lg�/�b�M�}�n��&���Ĭ2#��~D|�K�[��.]}�f[>f���h�`��$���l/��$v�(A������a$}ef0f�Mo������X�ZõM�����[����u:g7nS[�s�8���Pa�`bu�#�Zc�Y�/�Gǔ�Ɵ;�Bf�$?�^�&�i�_{�+��(0�^����ς�l�;�/�����	Wp������U��r�����c�~Q	�⮋/c_�$����&����j��*��2�=��*5?�6�F�k;#��|�X�Ş7��_J%[#�6D�ra�h�op�<eƞ�[�.,�-��g�6��E|��U[��V/+ W�'"�'�Axi[:n�/2|y�ӭ�w�vD�T2�e06GLW�k>�.�K1�cɑ����j��m��D�b�v�Bl���D�;�W)�/�1j[�~K����!�!IB�MU�>���v��QW�ź�mV���G��Fln�cƳIp���ϰJDmM�N,t~TӮ�;7�c�`�.�J�4|z���wJ���,�N�z1�wqW��UI�<7�N�iR.�Zn�`�un����œ]^>�/ <���ӺJ�������c5^-^&�i�=p���XL9D�`��J��yH)~�0�%��/~�'2�b�<{�b��l��}J��]�t,�bF!��zz�~z�S-y�ۚ��}���r��7Q�����68��Ġx����D.xA���a��oف�WhI.��e��)�#��W��y�6W���g�#�o��ӌ�zС3�}���A�K>�iﯬO�L�'5#6؄8��Bo5+�P�	|j���nYM�o;�
^R��.Wm��DD��.��FE�V��_�x(O�5�Y��_>.8E�]�_�]b�۹��6����2�69ؔ�-5���R3��RP��g�unF�)��ط\p[���s�Uu���f�#"[���le���,��Ў�<��Ա�1ؤ�{J� l�y� �|_i=P��݉������	U�zV{��'�����f��s}���@�V�����f�[�Ec�c�A<G��Z,�G'�/�d�c����fp���b�8M��jZ�j&Y�J�M��Ȣ�>>��ٿ�Xm���K��9/��]�g9��3�4vt�o0�m��W���������W}{�N�/N����TZ�f'���6t� ������b�/��52U�i�B��0?�!���R��S���" 55�5ӌ(�I�H�
���R7�p%�{�jׯ!Q�f+[�C��j�NK<�]�SoЂ����H�����6����*�`_�Q?����u-��|����1�̄E��X��Nj	�r��$�"�N�$������F:*t6uV������Ѷ����*맵�>�O	��B`��+�j_����Qcs����s���UIG�5���x%��Ls~�[�aL�4z��fb��,�|Ȳ/�g�f�R�里C��!O��%M7��� k�՟��S�դ$�w{�'�t4��;���I����Y/0�֬6l����}�QB��:-4	]��;�W�4�Is�]�Yg��$R���ExG<�kM7g����5��P�4���m���o/������:�ȎUN@D�_Vi3P(W�#�}��l���xG��	��{���?�����QA����+��c���g~%�[��n	��ge�����B�Λ��SA��AG\ѕ�%����c@�X�q�ޱ�N�
�\��{!��Lۦ�:5�;�7�!��{,҃�Ϋ}��s���N�-M�	�nbtl>u��[�i�B,�Vl��X:0�������>��P��i_^�K4s��EF6Z� AY�)��6u`e?hk��؂�M��ߵ �qf��Fuj3�����LF'_a�Y��]�����%�� �wCX'��ɳU3㹁ƙ�c;�=\�+܀�IR"��b������Z���]�5���6o5a?_b���Y�=W�z�'I7(_|��>�\Z�uT�l	w�~��y�z"��rݺi�@�DK�=���f��-���]M��uQ9'�M.��z8	�P�?��8 ���iu�'1�|&;;Zt����u����'ђ��7�*y?�OBH�>�m��粋���7j��*�L���A���ʀO�~!wZ��*H���D~T�f������%�ڊ���̥��Q�9(���^MT4���<�'?��y9�.��(�h��f���RI�-�]�a��
5[�����5�^�H��}q��Xcv��u�#���h�"t�{���!�b�H,�F�����y��"e��3���Vt�;P�o��q.��eE�J����C���V}o)�w�gzJ<꽸E+j� ��2�;��=	y��6���.���)��S��.����o���>[�wH��R�L&u�;}�⬢G����n_m�+�o%a�?�@%Ψ��1�p�|���ݐK��z��as��]6-�>I$Ha��y�	�9�;˔�ؕ
�Q��0A�l�_P�NlqU[v�c�E�_��+(�	RD#	 �gM�&����'�04��f<x��Eջ��L� �@{s��F����U�[{[�/E���{�_�A	]�E��*���Zl�*h�_�Z��l.#��1	�v=�����L��Aoj�R�Z�v�ǵ�ƫ�IL�����n�\���:�w	�q�Ԃ���k��R�M�����=!�{l7G~ϛ=��=��H
σE�	���s�������+j�k"<��;��i'��)�KD{�*�����rJ�_�����Ե����׵`��P[=���݅��d����z��Ô,��m���Y�'����M�����35���T&>�d_�
F��lS������P����K�ؖ���Ea�}�5
��H���G�+����l�?}��D����J&��Y��&6m���N�R9��v�bp��pW�'�{3�8 �n&d]EZ�I;_)��ܚ[���:�P]�����r��'P#`�i��.�o���e�Ķ�+�qHW!(�6���ɬ�ԅ�\,IU-��B��T�Dp�âưG��`¨}�E�AC���)����§�WI}xZI� l<Lw8���ݹ�b,,��Di�.�,&�i�z=��ǔ�������a8}=d:Ki�ZԸ��,T�@-=�껷CETR@tC�ϸV(�Nl��X� ����J.�M�J��M���V:�F�U���>J>O��7 �fv��n���ۼXc��QU��tK��G_M�}��q�;f�<��:��G=�7�C.��}57t��+٨5�%ȶ���t�� +I�q-�:B-DIOl�D�-�JH��_��ֳ�iϛ^*PM%����	v{X4�[m?��u�@eb#�@s,tYq��%�	"��~�
'v���G]c�79�����Ye,)�t���SA�!���{���jnt>�aE��0�[�m��Y_�&H2!â�q �A�e�2yqN����j�@���pz�)h�z�|xA�L�<�7�L���J`���6_����*`�|��^�0���V�B�(����R^�Sv<g�T<|Z��$#*�D��5ȫ��d:_�+�s-��Ъνzj	�v�[ى�9�����HC��&ݹu!���5o9�e]Xu�O��3�Jb�k��6�a�F~ �
]�Vr�K���^]/��@_���kg��N�+�ZN�L]�&��/�C+F	�QX���G|}�&R����B �eP��b��T.Ŋ�˼�����1�U���8tҠ���M��^��S����rJ
�:�[������K���*�vZ}HW���ٔ߄���(6�y ��t�ɰ�=��nA����X�찪64�u�J'��.�N-)�$�>��Goj�;�AL3W���0���OS6� �<Z�%�އ�t���H���I�v,f�
���Y䬨�@�>�@�;��^�>K��+�k%z	J����2�����o�.�O�A;�T�+<����>�*���9~���f9JI�+���Tdn�1��8�8��)�~����囁�Qp���̙�ʛ�y�ݗq��4��i�na,wgJ��e98�ݯ�'�5���6��A��P��
1,�� �G��|�ǀ�M�+���@��9#@;��Aw�d/V��g��~L"����0H���2�bq`�o�/�q�:�^;ϧ,���ړ}�?����}S���a9�<͜��n_��ܓɝ�ñ�M�
��V1ߛ��3�Q�}W؄�4������b�MS7�!41��Ġssg#���Y�UɜPE#^v
�p &a��LI߷\�E>vݚb��5r�$nz�E��8��x����1V� 3@�B����#���[���5��J?����k}�4�L��� 6B;D�������.���[u�,iL��b��h��('o�Φ71�\>Y߰_wI���u�7�"v̠L�&ݦ:�j;��)�<c����Hfm�}�2$�q@�&�x���ɶ�5%!���8�pڞ�Ap�"i-��!�Xg<�ml5a�e�}a��#��|=@ /��㒬G;�LS��Vuu���G�lC��V(q�
�#� ���ώ�l��==��xdoî���KY��������}�?�B�G�DF&s��~f���4�:%hY䓚�!�h��O�r1v��Lo�T�򟋐2Fr��K��.k�w� %UWx%Ĭt6��+[}��R$�:3���0j�i�g7��^�'��9?��Y��Z�&���e�灥9�t\6� Δ����7� �����[�p�L��	���y<QU\�c�$:�j��D�ji&٦1x��'h�'��)�,Q����_&����(�Z�D4�
�e�}��5$�-.m��a�8�c�ײ�_ �
JU6N�~��M��y�g'I?]%+ o�����=G)�t�Ν��l:z�|Xθ(=僭W���|��E)rXa�E!C�,D�E]fwĂ��ֶ�Q�-����@�JG��qa�<�%�W�A<��'(����	~���R�"��%��Hᛝ�U�H�zf����r/��5c�縘ܵ�i�am�^!�֖!��3�#�ąt�ޢ��%1F�_`p�yR�.�M�
M��#B��]0��+pl,�#��Y��E4��|���K�P�Q���V����PV}8��؝�S�DN����@w���8�I/D��A[3�.�LZD�T�܆/�J���52��v'㲖}E�i�.8�bjڹ�?�oh��kW7�KF]�Ȳ�[8��v�b�W�������wdٚ��{�Α�l�����UN�Ę$�0��({�(Q`��'�)�y�:�R�q�	3�"-��*��	j[����<+�)a-�.8բ|p �ɾ�[��$�z�����nY]-qO(ز�n����R��@#��rF���w(k��j�?�:�z�B�S$kCB��̪�Q�P..��%2�)�ĕL����p