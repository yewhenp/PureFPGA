��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ������Y�^ץ|Ue��1�*d YC�����v���7�/�P/>|�yXdv�֡�_F�6��tU��|#�&�!,\�t>���۪GBn:0�#ċ��|��m���f1m�`��fy�e�+A2�T>Wc�e�*�ʸ��\]<�UI�5voN����+c�����)Ũ
x*i��+��<����a��e��{Ekx�����lӇ�ÉϱV��R���ԧr�a	�_�2�UB�8�I �b�����K�m�˖��r�67���6g�T����zP<x0�ؤ�;�K��]��^P���C>�[xI��3؊�#�=�{ � y�����ٛհuzKȹ���r��빕��Vᶪ�{|sZ�na�hbd �����r��Y�rMP:��o#7M�{�>YI,mw���za���y�&:���zO�5�Ԗ4��p������Z���u�\�h�7m9�tⲟZ�lϽ	�y�-�����@ޔ�m�6����~����z!�7۶O�sy(�D�I�����L��m~.5�ƁE/�,e/�#%Ҝȗ��� 3s��h��ʞ�)8a������Q�_R�Ս���)��:�}��x$	�E�iPq�l�d*�.��K�זy���N=���>�<�� �H��*{�G��oIt��+��:w�2�=�՝�ҍ�;vm�!.V�ܔ�;�w�vU"���=B#��lt�C�ja���#R��.�qv�ؒp����S�7�ξ�w=�y��1�yEq�C�;��D��/���Ғ����k:ە�'j�/�?���11F��(na����k�q���x{�s��;���W<�W��Q��u�h��	}M�ʻ�����5���-R��)���B)���n���XGҍ��mJg_Pz��t�>�^@�><zX@F"�P�G�Z���aw,�d��^'Þ]w
Im߅Vo}ʰ��E���ɝUu��
��,�0�@��j�kD��f4���\��B��vmPx
v��x�k]�Z��[C*٣�|��;
�;��.�J�"�D���1z�T�p�s��#g��h3l�e肖����\B5zi�W�?����%�i�R��B ̆
�a���N�`�H���B��O�����O��ԀI$��)H
�ۋāa�Oh��;�-�ryW�#|�_Կ�)*���*��d�{*�'��J.��\~�D�n�q�k%������ۜ����"�q��S�Di�?���n�Wj]����OQ�eE�� ��t�{H����bq�?�s�dy�1��Fv#�3Pj�U����KqN�AW6�Rn��Wr�vC�;����<R�	�O3MP��4�p��􄧞o�b��G�)_FL���U��2�l�Q����9�V]�����O����>_���`3��@[Ö�E���F�A;-���VZ��\��P2�^��M/�T����r��\��᥆.�1�(���9s2L`�?�fB�K��>�)�wtB9�Ū�*���*W��qWN��? ���`\�;ʁ8�9���bK�X[��D&ī �j��A�%�\cҫzNf���"�S��W�3�I�Ke�\t����#8I�UV^I޳&���Tj���ep�	���3���9Ю����~sh��K�����9{���A���9��I�Edx@]}��~�*5�Q8�(�`�4�µ��H�1`k],�,ev��[/��Xg��zw��'�P@�s?pJ8EF�lc;��(فصB�˜�6�]�B%)E!��n����I&*3�*�4[�������g��tQ�ٍ�R�h���D�6�� ��Z�&:���#T�T���?�u��� ��<��G�vnCdU���P	���3-�P#���I ��!+�C�H��Q$�ٗ��}��u�U�9���ɂ7��,^czX�_a�*�j��-h�$�����]�����P��ޗCf� �����=Fc���iYn2�+����5P~���3�.�TT�{��i�����/QhyB�A��4s37!O3�����_������I���4��Ǐ`�Ҁ�۽pVz.M�/��^U<��V�a0��%�r���<5_#V�` �z�'�OŷG6��:�"m��ʉd.�Xi�|�ד�T��U���Wt*����|UZ�$���쉟{�u���rm�5�yn�n�!�M��l�8�@
VE�h#��� ���4@��9��<C��X��u�4G��c����;��+2+e�����![z�͓t���J7:6�)����\R�L
��G��N�q�Z�JU��2��.������ᔽ�ow��'c���<�!����4���/M�W�#SGnP�_ K�ct>q�/&&�i���]��j@�@��R앫32=�,��G8}Y'4 �Ӛ�B�|��?�Q��$����ņ�\{��E=I&��.�Lc�Q?�ɣ��Ti����B�*���
9�$���!�q�6�bAE�ָ�H��8G��	���<���_�-�y���X�	s��B�� ��1zeR��<���<G�VX9�&a;T�x����������ޭ�ם�޸�C8<MyX3*��f�����R�~J��ִ֒& 2F���E�6�E�_�m����Ɩ<1e-n�6	�'-��,�0�Q�b�}�/G�΀��-��oa 4q0`N�|��.��t�p6|z��4���at��h�D�T�X��ۘ}���k��u>F��S�a!�d f�I��N屹vM��h�R��Q[Y�.�/�6�6X�7��0M`�1����K�d ��FБ��
�3�h͊���P�� FY+X<
q�_��W���Vk�Ko��5�l��(��d����t��R���-����䜶Y1�K�X���
 �%ؙ�'����A��\���<Q�
X;�1��}DB�6 ܗH��k�w�2ɀ2�Q�A���g����+MSI�"�li#+_��Y��+�Ó?�e�*�(g�R�N��ۧ1��w	.2� ��鑞Wz��8���-۲r���̹@"����=�b�ւS4�4o"�##J����L_�/��/3�/���b�A�Z�?%곌�V�O��EfpMD�t��ү�p�)���u�Y��r��}�m�\���˱5���[��:�_�v{�hk�@��]���$j��8~�\g^�.��tQv3�})�SE��6먓t��!�A8y
��h�Q��]��������]�Ͼ�w ���C�aǹ՚��-�L�C zT��B-��R�=��5q&ܓ�E�&�!�`ٽ�R�2�V���7���^f�{������ؕ�=�:puj�|��1߅�sYw���x�(�ߚѳ�u(�U𨠼�F*}i�,�"��?b'c<p^m{��K ��#�7`�����#�-��u�01!|C^˨��]rA-1Cv�LxI�s��I�ʚ���R�'�I�)|��`WJ@��Ê�9��*
 AX�r�wv�G�
��j;ۤ�6D�&�\!hmNZ�5$��e��hE�v[�2��+��[G����#��d���H8-����l����ӂeM
���M��*�!���O�u�@��B��s��U1ݗ��P��d�KT'�xt�J�'�E��(k�e&� �[N�v"8��7�_3菅ױ^�	9��n��h��$�5J��QPa>Fg�~�:�x���U�#�?�.y�iOI��,H�Ho��m����F�S��@6׋Q�xwy��*HB����O�4�c"��u�.�L�����`���u͇#�d̃z�0O.���Â��/�s���9�+�1�	���Q[�!�ΙȌL��sl*��	M����K�gwg5B,��l��JrS�vAJ��.���x"�2��������'P;"�����"��|~t��4��4=�S/;����t�[T��pM�}{7l�4�2��R��[���>�1� x [Jc���[���Ȅ{S7��Pr�^�C�U�V:Z`{m�p�Z��F�9�>ۼ��h�i0��"�t�s���tki3.S�R�
��a�Mz���WV=���L"��/r��q �Q�3������ 灳˼9�K?�jI��I�z��	�K�\&��U��`rS�j����\o~?��v�)��&�P�T��?Y�Fm���>�%{ݴ����d-�L".�V�������D�f�˷����qM��6똒��ΪwXJ����'�uz��KB�6pM}�,%����oM96\��p�4@��I�H�_P=�O�>�Aڕ�I7�5�Pes+����fZ��8��<E��$x���F�6rxҽ��1�(,�&'�H�r�J�
�J�g,�/>	�u��w�gg1	4�X0���M:2�:!��~3�Ȇ5� Eei+ֹ��
������*�3w<v�K��b�克�����������54�#m��i�	E�7�;͉ý���_�Q�xo&P�I���Ob�+u"�W��@�g�Ӌ�(���̲OB�m��[\.,'�̹�P��ʃ�%�8k�]E�_4�	DjnK#thG�Gj�.�j9J�����t}l�}
]��J���U�'���M7���thsFY��(A�����8b�R���ɔ���P��sR�6��J�C�d��h9�Mv,���f�q��w��ѥ���	V�v%�B�����l�rv���~/@��I�Q�3� �u�6�]����X�?��]�9�j$�<�<����9#&�]�3�\7��X�4pl�-����Kw�9�$�K9�fS�� ��B���JN��2FY���)� k��Sɍ�;yf�C"G�nTnv�1�9r�^ii�ײ�RI���6���|�����Ƌ7��_~����N䢗�: �|_�)�^*��`����<��lr����Ga��f\#�! B='�5�":@>��>zތ�����]����u�دDoY��0��c����P��~�x:�P��"�*���x]x�C�m��P��U�UU=7N&�y�!i]���P,o���{����"��(�x�^=���k��M�tM�\H?���Df���\��4z|:<�M�oo�I�TC/x��'��+&�/���V��3oBN���)<��j8���������H�<�ت)�Y8�����T��[Pt�p����}��e�5�Bi�HZ-y�������'j�Q< ��:Np�9n�~9�������Q��g�|��յ�V%��*tuٰ�r�F/�|gf����k�lA�wkmm,�B���7>�J>.P?AY�Ԏ[٫�R�{	{Xu�(0���ȱ�m�?�o�S�ӰzW+��o���Nt`��� �"��4��K��D�[��c�ݺ��A����C6�4'��N��Y`����Ƽ�o3gj}�>M,.�l�Z�ypya�����X�_�y���&Lv��r�D�ޗg������i��_��Ў}�֔g�4c�8=ø3Ժh�
�I�T�!d���v��J���k�D����{���#�����R%$��J�>F�֒)�B1�ž�8�&◷�k�?�rZ�f��4��F�fKL�z0����6�#���
��V�"^��J�H�k[�OΪ��*>�#[s��+Z�4CV
�y(�
������.��-5\��K�{�7U3vp���r'���f�At݁51�v{�'�M����=������a�*�,���X�?c��_�!�����R��0�--�������^��C�	8�8��Z���m�&Hs3����Lx�,����(���E3��{�y�xl�6g& Ahʝ1Ǎ��+M���W!n�����ov���0d"���Y!1�:����E ���~%��/��,��_�=�������%s���PИC(���t��ܠk�!���l�>q�UB�SD���ځ
D�6o�����If� 2%�����p�����k8����{�T�ҍ� 1���?��`�	�����~�u6jQ��`����s�XdA �������+)��d͓�.;����чu��/O:`�yc�HK�ꠍ��t]�ģ�]�p���5�+0ha�T�}�6������e��8F��%w]ʟ9��e7�ʗ�3X��=- ���#
��������;���.,�Z�����o&��Ȓ�<���G��g�3���DV��l��4׹�ڇ��)�n�s�t
��=�ex�mɢ���N����8�¡>q�|XV.�i ����Og�B��b�p�����;x���P�i��EL"0I�j7��S��3��E��n�c�XM&��q���QK��j��N���Cr_G �P�e�CtTÈ�����9��bLi���<��s��q�7��4��>7׋7�5�/Й���̋��9��_u�I!��1������9:�;^;l��L�4��Jc�/A`����3�X�,��\�NE����SwP��F�D]~�S� -�X�&����sg�w�\�Le�~U������	�G�����2�A��P38����ߓU�8ѸS>�X���OsS�(�bYkR���6D$	��Tu�?g��X���ٕ�6?�!�wYWlF�ô��m���W�Lv7u�
h�%�V�g߅�8�@o�r��,}>��TO:��;�/旀�ȡ��_NU�؟V��N��eDs�onyW����ڱ�s�	�9�T�8y��F5w���%��!1�.](���Q{���h��qd�H����%���hfV��Ro�9ފ�nK;!��Y�
�p��\A�Hs����cz5����'bl��v�<�M���D]��oѵ�
j>�J�:W�h�upA�#�>���L��\#u7*��0�]��ió.!��{g�iF�٭��\�� ��v��o�婋�>5�ޅ6��Y��2���]�Vn�����6@Õ�L{����2��T':�J6!5�i��Yc��O#<1���]���[4Q���������N�%�Ն�����i�.+�����BӼ���Ǘ�X_ܞZu���=�G�k���q=�)�)����p4��6ǔ�X��Y�\�#^:/����>�M�&t�����z�ֳ�]D@���yT�����V?�
WrpU-`S��v|��q,��5~�*f��I��+H�}�܏@����2��%��rH�DGU�Jͫ(@�<���>���\�ř�m�C����ro�"�/��/���P�>!=F����t���
�j$��K%����lW��dX4+m���i��I�-��8�����5�E;X��G	V'�(oV�f�dC��޳�??��58Y��͓������܃����>,>��M��R4dj
c�B��5$}q�;�3���G҆�gNYE�����������BO�yW�"�Zx� (l3��:�h��(e�X .�Ma�p��O�eֻ�䈞�T���iTyk��*����u2�X��r//ftB���I'��<@=�>���&��Ϯe�:Jy��yx�T��Q��,�4£�8.]d$��\�Y�"ښ���1����&���/���z�=����hD����˽���������2��`-�5�8�;�ڃy�o԰}�֩0���!��C�3E�!_vۊ�3�6��]�k����N5Cdqѥ�I ��_�nQ�0罚F3��|3�'��/2>���9}�S��m��7�ZD����+�h�jT�6���@p�N�R�_<��Ș����>��;��1�4��Ќ�ƈ?���}|����V��wx��󎷔�[�o����'o�Tuz�m�sGx;\�K���I+jEL!�'QPq�����+.i:�=9�,���f��V�4�j�'M��J��Qyzᶚ�p/z�l�w{4��eE�'��ۯg��9ގpJ���43ٴ�Z�q{ZZ
�aU(��=�<*3J���P{����L�Z�$B�Y�◒��pS�8�a��<2�!80���ՙ��\"ȽP��d�bm�-��g[�
��v�0�娵����>�z��$`�@vzSmOz!�R�l����3-4��@N:�ݼ�*�HY�s����$HW�!�(eU^�n��
�
�1��B���k�r���ajr�<n�p�ʃ�ώ~�"	���~vO�c�b�c��+��b��*���<��0�L_�dc��L,����#��#�1�C�n[��;v<^7Qwܤ\	�5(ͫwKȥUI1J���+��׬q�V:�i$	f�x�)$#�.�b�BfqY�
x!ݎ���[���K4y��dв`�Ʀ�>������������P�'K|ue���.uI]ByA&�����j���÷�(�m��zL�*�4��]���>�M=��}7�g/�Ba�Ʌ�MM�En�r��=W�YZ�1}��w���л7�Xyf�n��l�|xe5K�?U$C#��Z�f�K�5�L7��k��a���9��ȿ�ԬZ(�#�Y��|�&�Xػ�u�=��ҚR�kL��I ir�f�	��L���B���-�6�h�8 ΐ�𖸳�	Ӧ]�x���f��9H!(!@�<���M���؊�|(<U�����~�����si�p�H�A��_oo���w���@0\�m	���%�ް-炢��I:���F1)z���JS����|�$���#�{��I���@����n�쳥h%�&eP ��Õ7�9����^#��j-�py2~f��Y�\�'���=we͵�ܨ��E������C�P�;�Ȇ���B�Ԟޝ^�1t�Kg��ѝkE�;s��Vn�V��K�qx�+\��`	W��bo��R���]Wy�o��q�H��U����@�T�\�e�����"	�����*4j26�!����|��%	L�!�zy.����ak+uE�]Ѩ�6�@ET�����h�Qn� �R������֩�9क0�Lom���88�s�.
hY*^��έI�z�k�US�Ox��%g�Q�_��ZOЛ_����L������կw������Dǥ@�:k ����i�����	��g���I~�>[(ĩ� 
r�c����pD�Y*8X��ӸV��oǇR
 {��}5��@oV6�ŜW��	���q͎�����B��2YG򢡑
����c���&�D�'x��I�p���m[�\3�.�;��hV�[qc�?�t�ýg�Q�U�J���n���A����c%xUL+��z����5^Z� ���8-��R2^��	%����%vq�V���'�rT ������הRM�N�y�jq6R�,������:�!���rX�?q%�]/��>w������rY�j�;);gt )3G졽;��H���b��'i���.�#����{Ov����{���s{{�}!�P��8q�@>�H�eI+!<J�Ǵ{�m�ݪ�3S]�/Ҙ�{++�і�'z�Gz��ޞ�V�ٗ�U��,+&K��50�arn��v���ϸ���@��C�+������8�n