��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ���\::��_5x'��n����%N�+�t����	q1��6�1b;��}��Z��>8	z����6t�Ө=��͠v]C	wi1�s5i�-�iwi�j��|Oe�O��T`yI�R�����E{!wva��o�����r`��5ȕ�L5��^F?���q,�tǩsA����79�Es�^��m\�rL�!o1��is���+@N�)����8���L�Nq�C��p�}�P@�� ؤճ�jm���R&��9RI�e�Sz�o9d\Oue%=n��npM�;���}�<�ܵ�!�N͆����?���t���_ܾ˯x6�x��%ұ���7��8T�]���n+�oW�~�_S}�&AV98�|�瘵i�"��}0��}>�u�i@�@T�c=UQ����xIV�Ӳ��p�v�&�u����6?�T7gy��zb\��rج_�%�f��t���: )�FE�8Xp��E��1�*��'�Q���1����)U�C!ZO2Z6���ۤh^-�	�����?�b��b�#���{X�eUᔦI�R5^�%��5N�����F��f�J�ќ�	��鬶�s̼���@G��,v���Py�7�O���yIQ�[~X)@��΀u���4��ǹ�z`��d�g�Y>���d�s�߂�}6R�]*�P\N�MY ��Eiq`��I�,�3a��ԛ�H��K���|�*�.�n���4���=��\\ �l�9�b+�<�����e�2j�	�L"{�ͣ���߼��)&����U$=���z�����U��I�q�#ģCg������Nx!�4�С��6�l����N�`�� Wg�	k� &d@�C�V���z"o��kO��QD0	C�E�p�N�혃��Ŭ"a�m(�wb�w^6�egj��f������v�j�?��m+���&6�!Ŀm�'�֣E�n�����ęq�!ĺ�e陙���HI��hQ�Fa�_�����'�FZ�c�/ll�u�z9Ǽ�_�O:�>����:����ն�,3
����~3M�a�^��]�5fN7<q���kfG�٤��i'c\Τ|���=�#��^��fFΊ�;�]`9迎����hO_��y��р��M/�ٮzw.vjF]7|����
vWUcëZf*U}ɸ����W |�#-��]���ںh�����6�U�
����S.�?#q����5�#xn��o@	��>s�*
W�-r(��׻�.��ύ���y7�����^���z�^
�6��һ�Ӭ׷���沇3��v�ez��57I����J2e=W#{g���C��>[S����1o�aV
�����@4��8_�׉o8�tsm����J�ͩHq�C�QFM�'�$Z�Ц�f��<	�On��{bu���?­Qu}'�p�"���8x���W7�/��o�S�����B���-QTU :�g=�4�5쥵F�|��z11Yp7�$E�du�@�H*nz����D �ϊ� 9�5�g%�h�0��y���������ğq�%������_$JY�i�j�^�h5�|�)�?�MU��M����}��s���Kv:�}wk�d]u�F5�O@�D�M*�8t�I�r���q�H����['٫�
�(X��>q��츺x�e"�aD����<�ǉ ���oGP_�ZC1A!�s$���|�n�:����{H�d�����Ď�w���ɂ6.X���;J�1�%L����&�ԅ8](���+FM�*�"5��$cN�����Y> N�} �P��Ϳi%|��1@t���K��ϖۮo�^�"�l�i{+��EwI�L��e�&���������dα�!����	]�*��!�k�Jv/b�0�+B)��]��}���~�ѡ�w�gL_��}���{jOZ��y�d(���F�TGnh6z�J�+Ld����&k)G�v�=N�"b<aI��C�6dzU��iu,X�IZݛ����h���5��֘�I�����������u�L̠���6���J#�ؠ^�A�w��T���r;;�^�?��������(��R���j��x�{�|)P��c�b����1�����,=�H���M�o-�SX3�����6.L
7�����q�l,I		LR�!0^��Q�Vș�t��M�Z���A�(.�S�P��@�|k�x���X�I_�|]���=�G�a��td�y��4��DW��Ҩ���K�$�R+'��߹�����笌���kM��s�n��!�� q���,����wd�O�ؾ��>a��	�������y�uY�w��~����c���q����A� ��$B-d���G�>��ܔ�ġ7��$����F(�/�4s��٫�3-W�M,Q�����Qlt+:7���_lT�8�	�6
#��Ёb�����R��D����X� *�ֽ���qc'x�\<���g�q�)�����ۭ�2WǫY��&���X6��v�6o��|=Í�F�Gi���_���̓ߖm�E��Km�B��3� �4�y��p"|V����PA���G˸��@��@�iLȳjb�4@Ð���b��঎`�O����#f��U�-��'qȢ��s�~?�5�C�+�_��Ғ���N6�@�ЈV(���1fR��z�0������rp7�=�E�R6������S�Wq��
Q$�ŀ�D�n
_�4�O�����۩f$� <�e�����Fx�¸:F��p*W�?z�Q�^
#�|��F5��sЭ�"j���)JoIn�A��Z!�<��8.Q�#$��I��{s�D��I�ơ�1l�ڊ�xxV�a��gc����!cS�Q�6��Kؑ�|���L��#Y%�$o�B���:>?���yKk��?�'��CZ�����(��Ր�9�Н�<�5Y���;}�8�!o��ԷH�j��Ưg�c����'��R#�� r�amI�Ʌ/\)��j���A����WOΔ+��3ƍ��8�V���D\�;ӫ�+��T�I���b)��꫖`W����.���e#�������?�d�&�2|d�]Ƃ��� 7B�s@;ʩ���4@ABS��1x��"��)k��X��tz`)�{-�8����_\>��t�J�p�h=���t /D�4(�-���Gdp�b�<�kf�COLvԊ�u�}f@���ab{3
�T��P�p����m@��yd�.)��L4� -�o�A����%Z��Ġl��0-('�T�����u�Z7�B�D�P*D��F{�Ǜ*���3�d���C�����Dά{y`�"ʂlTO��g�8�xb��ڂ�|+ߴ�L�HK1��>���ϒƣS�|����x���E��u�w�L~ҜQ=��d���=
)uM��:$Ӏ|R��A`�~B��K��xr�u�^uqO�Z�h	��a=<�9E��f��z�f��
u�,9���Ӌ�$l>'!�	M��������"���rc��k~������������ЏMk�,_*i���s��j���A�/3�*�銆+0��
b3g@k��i��D_�0N�M�~�*�U(D���-����9%B�s^�Y��ʸx��|6���~���b9��1.H�,�T{�'�����?���v��,&��vtM�����=���WG2OFЫa�����^ �K�jnH���l���~�Mv��oL�d�b_����:?K�KԘ��o���3���zӏ�0��'�G��rHB���Mf���OF��l���y���))��Y�a���1�4�ln�)!бh�)NLYR��#߼ѫ��٨2�C�aLV_@������b9���Y&ߊ������6 Z	��\�f�{�@��$�{�,A���4l���KG�Dj���_�q)I�w��'�k�}vX�����ƿ� �`8�5�<�8�x�����*�tF��5~�<�y���!կX��j;�G�"���;CQ��h?%�W���O�XY
T�@��^�/��ԉw>���42b���}H9��3�>+(�hZ��d>@�,�Z��I^tb�GRB�u�FS'�zh��($�`u�����;��~���-���W��ċ+�48�,�Z�'�(���
�tL;�.y�Ѿ��X�kJ�X�Z2�m������h2i�#Y.L{�K�w�2�@V~�ʂnL�j��8���������gjN]x�mhC���(,��6"@�B�m?���2?t��1��[rᑟ���ٻr�c�u*g�͛���r�nD�X�U�wgc�ã�s��(�yp���ܺ��/#�>�G�`�?�����,%B$�|��vB��@��S��6����rWV]�]I&z�tkB�c����<`��gA�`�l_1NS��Y�=D~i.�5�
��e��;nr����K~/u���T��KHV��-�g��Ԁj���CNr>�g	��n���.���h���iq�$!����@|��٧K/�`��5y��wyN���������q]@eU��绨�Z~����E�'���lAx������Y�P���¨"�Xo�*��Vk�2��&��-�?�'�5#���8~�
��`�O%�ʤȚ��'����ѵ��)���2a �H�
�)��Duܔ�t	A11�����}��Y��B�������^G�l<W������3��$�ǵ�t�v���b�͹ssg7S�U���Gqv�NH�]0-�F���i�OAl� ����6Mzg����k+LV�3V2D��9ksړ����H��!Z���w*�|C�S w훢����`�-mS�^�6NT0�y�۞��%�)'FV�\�왔��4X_A	��ڮ�A��ü��7�C��rP?K@j}�[�ZK���7g�CP��kʱ1j*��E���4�����\f�%���ԯI�T��ϝ�J_Z���,	օQb����P�F�Ĭ8��ǆ���%荣/]M�a^��Q W��*WG���]��{�hG�v�r�,�#~�^�������%Ǖ�Q�j�C9w���	qkz�.�q���HZ5b����9���|^藜
ߩ0?v�ҊH���t���vҿ��� ����$ �s�]���q}V�5��i���y�<���C��W������=�J�U��,A~@ґ�i�&YƳ�j�{F�*��W����_F��R}���K��<l��a{�.�a�������U6���#�Nu��*|�f/��c%e5�~��?�J8ɰ�H������J$q���>nd�L��S�fV�SGU>(���`�5{X�G��8��2f�e?��}J߳���� ��	�ѭ
=hq���E�w8a}���F���*��xۡS�x�<꽼��$��Ԯ�P�2h�V�m�`&`��pR��a�x�y���q�;�"�=��Z����?�J~���;�~8%x�EH;v�3q�}�U���3�w�E+�`[��XAc���ڵ
���^=�-Α� �()�3��ۅS���j<\� Sс?Q)[yh�gI
nat�ڿ<R�_ ��v�o-ؿ�����EE �.ŜУ�\e�Gz}K�(���y�BK���������+�$BT���m|~�}>�T�﫲?
!SG	ǵ�N���+�W㚡k�D��}�v�6U?k`텹枏�$Lc A4	��M�_"�u���G��~Q�a빯�!0�օ�h�m7Ť��Tç
P(A/�A�=s��r_����ں�گ��`DY�e���V-P��ƫO����� �
��Iҏj[�1�v.�� T ���� 1�|��
�[�J6�|�?��s�ƫ*ZI2:�sz+	#�@�%��vD��7�Nf6ԬT$��
)^��d��4&��x��mP�<�˸� ��ќK�8��Qv�-��:���}0bq�����]�WӐ�3dVho��B�Vq?b���u��Xo�,k�i*}�@oh<Hv�[��*ϐ�oQ���ra2�����~i~�����@�AdMu[аA��"TG�Bz�K< ��v�+�C���cm��S+� l�Wl��VB�#*��E�0�^��R�5�z�+|)�;�h#®�})s���s�~x�hkr�)-dAb�J�t;��2b�~!����3�Kg:��LNt�w.�<�>��,|�&aQ��z	k�!+��P��,MHI���O���?d��/K1���F�n�ߚ1T@�j�3�q��LҸ~��W��}��ZR�Ymx,B�e�����Ł�mOa:����1��;���NW�&^��y�A<��)��oT�zvo�xI��"�O��>W��{��,誷?X;Q$�w��&^x�N��H�i�g?�-Ap*�x��N�g^���Y���"A�
�̴�[���>�Hz�Xw"l����u<��'���.�o�'>9_B��.Q 
<i�1��P��~!�N�p�B(�"K������T��5;L�t�y8JyU�zH@��֧�-X��82�0
� �G_��`E��p
�Ig�0׬��~y�~���~���N!���Ϣ�tށ�w�z��:�&
��h&y�rx0����N�O��i�\�%4B��bN3�/?*3��`�Q�����{IÄ�_�v6�D˼-�ēa,�+�i�l���~�J�F���K/D��wd�f�iԟ��0��� j2ϻbF|�A�H)@�Q����rVK��wf�����CR��w8�>��:�/�G�ք�n���+G54�2�F$�E�q�6���Km���+Qm�j�ˢ���p��+ǂS��E�
�;o-�l��2��${M �`ܿA$�ċjW�����ָ
�Dj2���]%�����vQw���w\-;�K�}H�v����(��C��}��1�f����.ò�|��E+��+Ft�ʻh����2��%�;ֱ�!}��(%�;^��P9��Gk�z0[���a�2.�ʱQ��H<!�a���)�4/�5������)sk%r~���%��/�9NQ�� A��M�&`}p�?[1�׾��&�Q�r6�	��ƙaCT����e�=?<�S�@��������h9}�!�2�.A(��Y��2��Vk1zX޺����ˑ4��.��2� }��V��Rx&�ī�i�@��7+�5uP?W'�y��Gn��,5�r��!�777=�ӏܳm�~ �J%>�m9��+i�1o$��3D�u�̷~_�	2�n���7���)�M��y�����D��Jx�<��@7��l�yqǰճ�����iF��`6�y��3����U��{���8��/�S3JtK"2����������v;��[���4i�6�FH��V��b�>����vf���,S��n���S_AH�o���Txg�Ys�Q���J�}����FLP��ܮ������z��,��ԃ�(����f{�]2O�H+T܁���Xx*X0c��_,� u�0�q�mZ ��v�\�ЊM�Y�&�K)NIU��2L��|t�2�7E�����-)�wʥ,��aǲ��5�Jɾ`�ԾY�(OER�B}S��3�C``K]�=�D�-1�Hx����D�0]r^@�Ic=@�2�p]���L� W���;V�?�Bѩ3,����\[����\���q��(	��3!�t/i��6��y���O)��u�5���rk�?c��b�� 1�_�̜0KI$��^��CA#/�mJ�E�!�I�¥�0a�߇��ED��ձ"�ׄ���+5,�4��=TZ��+X��İ�/2>zۚCr�)
�����R]�~ �'>'tI�}������	z�4Q�db5u�`ɵ(V�K���L�D�s���s�Ve+�& j�ڭ�y�?$-��{I��W �� q*�eDQB?��a�JLy�Hn2x7DJ�[9�;�4/����\���PC�e!(�~��>�yFi�TYu35�n\%P������[6_��4��m`��"�f�b��V?V�dT�M� ���YmtU�y�m~�Yy�l�~Z$���+(	�/���9l�We;\���i^���L�s�2;b�N�9�bW"d���ѽ�5��*��/s��_�f�,�_=�QB�J=����)��9��.a�uk������d�/�M^���x�D��P#�PQ�������[q%$�q�A6��('�5R_5����ZT�L�A�d{���4����K��=��k��|�>�zs,�J�&ny�YM� P��Y��tyY㺈��)2d٠q��{��Rt�J���a�9[�^.�-q�83���5�� ��� ���j)��X�U:�&�gF���&����O�+�]2����E�!���A>�p��f��G�̶kI#��5�`�^��\L��mH�/|Y:[M�{�v~�=�����k��O��b��}�|�xi�&�Q-Ȇ�P��ߓ�#�<�J��92�}�i{5G&2ޗ�F�iZ$�_-�U�?����\T4;��96�~���ԉM������4a$:EUD����N�v�Zf�-2@8:���#j���C�Y�dI�艐(+�;fK�ۄ�h�De����7��xSR"K��ٛWت�:bݼ�.�'<�fO������>�-��7ľ�}nq~�)�0�ӓ&�},0]L����� �bxԠ���ȾZn����y�d�1Z�����z�m��hA��D{�����ʰ��ib`�\�;���B���!��I����;�kM9���ſ>��e�u��p�(y�����!'P��o��[h���;�e?V:L���Deo'���O?�l������p�(
�@a�#\��&#�$R���zӉûm�V�#�h�2<�TH��:'}�n&��F��������;��3F,�N!ס��r����������o���� 76
�7���Qe̖3>A��Q�p�|�@9�c��]J)o��xTa���^��%u���nb����I��
V�,,m�\�� G�[�P`��56~v��ˈac��֥J�ˑ d)c[`' ?�vx��g�E��:Duw$)��eM[��y�Ojb��
z&=<�I��w�F�hh�C��٩{�D���o)�����n�do'�:$:���/�Xb�u)�5�"�ԥ���Y�Lv�S\M3%��tk����A����Q��Ot��н��5���t�U��$������N\tUv���c�j���F	�����n;��q�0`(����#^g6(�0�[�ɩ���C��7Z<���C�a6.N��a�B����&�J� �8?�,dA-6�3L�����H֢��.9�#X��u��@4)��:{�R�C'%/b��E�.�rG��N��%>�~��<n{&u�������=��P5(��Ed�q#  ~�%
�"�˭�t��}�۫l,S �tIzH3�)�X��hSۢ�h���m���r��CU� �(�QP��+ŀs� �	�K'!E;�$��{S�Zp5��*%�I3��-�L��ځ��a)����hT:��r-a�f�X��w�3�(�(f��y����*�*]��U}�Dh���I�iܬr��ұ*G^��RO�/eW۳�hՉ������J�<��;G��7J?��g��^�����ya�7��cNo������~�E��� Ro%Ʒ%�ke�i��_o����L� M���WT,�V��UE�9�,���y�@�>�����L��4�J�Qp��R��X�h%��؂�<)HQ	�L�ײ�+V��7�7@���%�}�Q��Omv�A�.�W�&��g
V��s��pvR��&�߹�O}�O*qz���m����懹�&Y���H��t r��Kû�@��>�o�G�FN��8Y�%�a�M��,�� U�t��A8�����6o[����o�ߴ���ɹ4~�ؔ
/�	�Ƚw�3��l/��h��b��l��K�L0��UhgMΑ����da���.�??��2p)z
�i�m�M��(��XU�\p� Y�;&���}Z׽WCp�Wc�޽��b� �ٟ쫰��Q&E<�����W�����t�
F����E���TT�1!���#�oӿ� �Q����*���xF���j��tqߘ���uZ���6b�d��a���L Q��I�������x�^/Z�~��JP���S�=3N=M��1�Tz�kz�#��@ϸ8�����,��H��φ2p�;��ҳ��P�Su�-7�".k0��o���HO结�����*����[_��6��p0�����E��.<��S������8[�>W�.r�5��%��G� �Ė��
�Ժ���aZ|x:j�K���wO�ʋ��N<!{����+�y$4���̮�L��q`&��˝W��!I���L~�Sf�g�<l'���J*3/|��=��"��������e��Ǩ�.�K�L�U"US�b�����6�B�����
��F���Kh �c�R7����ɚ\"W�_��ҝ�{E�@\Sv�a��gm6�H��N�N�
��f%u�ו>߲�V�	�w��vkԒ���OS���v�����m�h��u���]��^��u�g�|�gx���;��ezb����Yу���Ww<�ӭ0D<�+1���7�&,���1$�L`�3X��
z���¥��{�±�)�9[m^��(&+�	Kg����~�_L����V�>���KZ�<��a���4I��0�y#4	��c"��J�ccd���;�ʰf�d���A�w$x �%^�+��������##�05���鷫0	��l$�XN%k��)8b��TN11���{��Jo�"#-怆DsD�;�_~�ɲR���!��7i�a) Q��ʢ=UM�� u�EY�P
ESF�ǿ���៊����*�D�J�d��n�����.9]�ʁ3�\�s�*uw��Wx�H�ƗZ�sp�0�ոǚ�^��q:��j�>�lѰ�����H��ŠM�f%��o ��FYp�!;��r��$�˄QX����g>i��߮_��0䯛�ʄ�4+*BA��ss`�k�4�!���:�֮�Y9�O3U�Z��R7iV�n�r�\Sŭ���"�H����TzO���D�h��X<��d�&.¹Q�I#���(=SX�vu)�B����c�s-�ƫB��׉9�[r ��*gb�r_����-�\Ib����h�T��Z�m^{Ѣ�\x3��3ŵ���M�-�RY`�;��u_q���VO�󠫶8h�7S2�y�^��� ��<�K5��� H�|2m����F�mI;V�d_��)��:ͽ������gm�6���)�B�� ��G;_7-2��1�G�̈́Y
y�|�Xs1�!O�Iw=N�*�ysT� 3!;�|�K8Ov�Ȁ(z~�6�N߸a�8�Kf"r��=�1�[S���
Q���`n)'	DC�&7�U	���+�&����S��h�^~ ��_�J!�@8xj�1^�=�BuJ�?���q)�5�
!ڔ�mZ�{��z���ʃ�[��PTDE9�R��0���bS��G��!�E?Sf�#B��M�Kj���&U\��V[�Zs�͹LS��[>����=,��:��	���
 �Ҩk�h�6ғY��8�ǡ	RbC\XT�U�F@�;$��?�>j����#�Yf׊hgI�`$�&�� ���ܡ�	2�'�����o�j]���m�6����[gF�D��5g�G	��W��ȇt��Do|�1'�d���`oN)���®��/HZ�H�H����+[ꄏ�N�O��S{���
asc&�|"`���d���x!k