��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� �R������JCgͨ"������"Wu.��z����Q��U�����������T��+Sq���w���1������*y�e����h���d���4�{:�ݟ�U#���9(w���߳��� �:ӱ�5�A-��O䘢X�,��2����Z�*�.��g}�T� �`��62��~�!{|O����ؔ$)�.���XM~��J�P���n�TH �E�_X�՟x�u%���ܢ���+��`فx6�<�0\�:rn�����p�!�o�}o����H����VyO�k�*�y���p�6�~\,��p��}B�t1Z�r��-�w�ҁ&�S�wY�G�;�;�)i�Q|�{��.u/���\��o�t�����Z�C��$F2��>��s���D��Έ=�ς����2�ʍa9��"�w���G�R�v���F��g�̂[s3��03��&6LƟ��5��$oD��k;�8��C�+�FE�����i�7����aZ��� +�f])��w�e��d��<�e�Y���J��E�C,���|_�T�ܞ;`oo����j����`� 2�|�d���	�l�M�F���*.�>�l>ǤY���֮ju�@����eVE�w���q>�2L/�y��؂YlW�G��%�0���m�FZB�*���#S�{g՞ z�V*���hL�U���u�L(�,�>�zb��+MUF�w��y΄#�P�w�*u��`i"�v!��h��h3%&VѼf�ɑ�L�_JM1L��W6a�M�i����)��l"n���&	h��3��ƃ�"f�*��޺+
�U3�Y�Y��1�nj��^A�}���D���a�k@�a���	����f���������$#��#��v/
?z�&�҈��=O<��r��j�2�N�ǹ���'��2�����x���pV�nŭ���/v���/��yrx��{�&�Hz7<a�P���v�1�y1$��������i]ލ�Z(!]���)֭(��2QvX17�j�i?F!%N�gZ�����̪��(G�g�&�#�RX�֎ܰ�������>�A�Cs`Eg�����!�:�]��'��4�z�(c�Z&6�%��a���#�%�Ff�4��0�sC�R��A��ħ@q�EUj<��Z~e�_�D�۝��LES��hdR�[ ҃�.~?�I:
��yƷ� R��n����y��!���?R�c���״�n��M�B����>���/ߠa�\��q�<؟��;zyy���@#vh�v�m�1��%(��6v�*���!W��Y=�#�7�Rr6�A`�.�(>�֤+S7R�^��p�֋���^�	W�EAx��gW�ܼ����H�h�@�H��;�Xڸ�j(r�U�M~Н���Vp��L@V&E�+���	Tښ�T9s��^-='0�#_�ەl�\}�¹��2�:<lW�U�����W�f�+e{��*M����e��_|o~�S�7����BŬ�0��f^��`{r7�8��X�wOr�4U|�H�è�l�,K�-n@8J�fO�Rs;�ڇ�Gx"��`����φ��:oC�cC?-�����W��K��]B�����Dϖ�o�y2�q�,K��ƺ}ꜯ2�3�������Tz��"L{-9t"�ǜ���q���w�k��F's�~�l��i�}RY����D�NBhL���ߌ�wDA������`X������~���^����v5�bd��/�3<��9�A� ��ɞ<��W�Jp/�|z'��݉��4דn�(7�~�n�~H������(�6~�����Q��ޚ<?[��J���Ta8�\��a3����"(���.j!��Ѕ`��&�1$W��.~Y	d��\��1T(��<:������_���I��{�\E��`۹���^D��~�5��n���g�Dc��B�2P�2^����`k�@�c3H��vOh�X������i;�2"��.�͏�K��yq�j8q&Q\��#�T%ѥn��H���_}#��@bS�:.ވ�H�OK���IX�8z( 8<��i�Fα'WP�e�)s�+O�Sqڎ�u�	g!�����&l@J�S�Y�M��q4_�n��l
���:~T���*��JOnu�)�L"�M�"�Wu%���듣A�+Z[D82YQ?����L��q<��<�֟�����(^�(��u�x�Dz⻥-��ʠ���V��)&����J��,�æ�-��*{��gݛ�hih#��\2{w��׸��9M$Je�W�_\"��>����i^D �Q�o���&���^bv�HK���N�ʺ�5\�ˤ{%���2}xF�q�����p��)� N\o���dPn�`bQ}<�a��V*m�(�w����*����0m��6BxP�Bc�^�|n�-N5}!Qa�����{qJ[)p홺�jTMx�֬��e�Ă����q}�k���Z�'c��"�����v�3(�-<�/�����
㱋�rݶ�����MA��,�*b��$t���Y����2b��p@��^�rE�@��x���Wb��h
f	t��3I�[NV	ߘR~m~=Jɝ��,�G��[ղ�
����I�y���_3�c5��|�A'����UE��d�@W詨�C��k���.m��V�V�W4��8�祽6��������^�51��B�E��A���M]ᬱ��FL���7�e�|�oOJr�GPLYN������S�
n�.´��d&���M�9�����N׽���K�]�t�I$�g�V�nQ�}$�Zʖ!NJx���m����H���w_�)A���c�֪�E��/�8��p9���|�D$%fi��(H)z,,:F��!e���f��4hF�_��N��Eq���Xml���x�.%�;o$�������Y�,f
7�����;	ɀ���F�lǋ6}��џ��"  /#,�-�>2M�*�T��h(XI�t�NH����
��UE@��5֖�4d�^��uv�_�~�^����܆���x5�{I��U�H���!�mf��̡���Ҧj`K������-��R.�^0tv"Ee�8��[�FF����i�r}k�۳-Jױw�!���e?�C����(�xn,���y�Ul`yA�HD�F����o�'�n*ɐI6-Y��nnx8�����	"�>�Ԏ��/��!eads�=�-�#ӈ�|(7]�]�u��ZpX]Zz���"V=�{�'�gY���� ���	hT��&�y���k#���#�S�UV4��2:s
LQo&��� ��+���KXpښ�6�6�P�#�9�$�6Ļ�N���#)�S�J�v�F$ef�K��j�l/�_7�ى��&�KL�D.���$�p�� �׾��Kяd�4'�)7~qȾ�̈��&{H�Wk��!��r&O��N��[j��]1gb
W8U�NՖٛ�Dˁ-��8�s.���h�v��as�;����#�(^�=L����� v	�����>��{�H6�,�h̸DŐ$fc���P�?��ی{2�vf����^Q�N��h[{X�y�Y�h�e�P�75�LǭJŢ�Ɏ���:��3�	�$2+���2�&�}0�?��%���m�4�U��:H�˛�_!8�|*)% X[e�z�
��-+g���8H2�RH�\'kG��+�f?F���+��͉����˙�1�UT��Hq�ַM+7�=\�!�B�ʇAL�J- ��9{�*u{e�����#���N�Z�]������sH|A+��ϼtX[\�'��>���'��y�U(���o��I�X�Ңfm���im�\Ma��D�*wá$ا`�n���r����4dq��LiJ��tx�}�� ��(��������r�����v�
c�Fw�Pӽ�~}��{I��%P�^���P@Xd]��2�s�O��	�D�*�G���BHk+��������D�S�5ق �A'�_��3J����ħ�I�t�f�O���3PG�E��x/+�e,�fȮ�5	����e�W���Q�-��_@j0Q����Z�ӤF��"s'R�"w��(��ܑa�Q)��Γ���e��%���@�Ȫ�?��H��^��9}�:'@����
�E���Z�P�P���wO�0�lU�[��|��V��%��˧g�$έ�<̤�)�:z{�����KUsK)�[������u���C6���s�
cC��m:9\����^|��X��w������31����qG�	[���&Sǡ�Ys���sjǚ\2��*8U@�fqһжاz�F#a��oTC~�~�(t0��'2
Vސh��,�pɌ�D�C�E�����9.շ�6/����n��ӱ�$���G�5�i��
���)�3P�u���5K�yq8Hp��f)�B�u��Mͤ��'}`VMu�!��O#g�8��vÆ�5[waN��P?o�2���k�I��n��U�"
أ�Z�ac�8���<��@"���w����`��}��O���K4�o&������u�`��K���RA<�7ȭ=��< �C܀�՟T�O�Ga��a�P�1��<�L�l�^,�
$^3la�`��@B\�fu�r�������P�Ǆ`�0�I�	b*A�"q�(�� s��p���D\�>��`�"�%{6h�u}�RҠo������z���+4������ztq0��m��˘�
6�Ȑ����vF-��	Ti�&�y�5;�jX����T�5i���G�wY�*�I?9u(A�lɸ�������`�;�9�1����FJ��>�d���ud�.`�x��p`O$y֟	�H�bN\b�޲��owd/)�9a$v�_��W����b��_C��v�u�R$���(�D�0��vDJ,F����++�`����*���~ꡖ_��� L}f�Ȅ���Zӎ' �M�Ȧ$���$f��t� ��km����h
� I������:��_����!.�_�3��}W*�d|K U|os]K)W+E��ܟ_]$i�3�PHg���7�b��e�%��
 �X���oM�I&���!%D����WOF�u�nZg�����I�B9�ͶTEO�� kB���h�r6#��΃>p��U�*��x�s�_]������Z���Qah� ��,�g������<$����2A��=��5+��v�L�c���T�e��0� �}_b� �uA�����,�btJN�Xa�xinh֨q�$I�0�yd�^|�5���(�z���K,��ͳ�$�HtO/�����E1��Ȏu��jI���׺s�1��&[gb�[)��2��^�����~�og���BIpݢ2uG��qd��.>�[���k무������<̽}��ظ��B�=ib��ᖏ�3�DكaP��i�@K�[��)+�5⋽��w��|E�� ��0�HG#��}��� �r�,�b܄3@/w�#B8���(��]�*V��/��(���ɍM�;c�'�௛Ta)r��[�׌�>���(��ue�����ǢcR:�R7�-��f�G�������Z�:�Y���� �y�8pQ�ga��^��v�B���K`�Bg�?-��!z�:�4�ѷ�M��J#���r	��?��H��m`�IO7x|O���#mJP�0ٞq����f+��)�����;�t����)�B�#o�ۀ��5{���X����q�TgK'9�D1�)�����p���bfB}N���-x��(4-_?����A�`�U�tm>i�̆<}YIٻ�Og ��nj���bMz�}6A�J�<�n+��+y&�t��w��T[�'���}xՈH��J�f���NW�lP����ksa��N�>�"��TU�L���(�������ߨo�����RT�t���#�ǧK�7����{�Q�N��Zh��h\�{%���1 l�5|U��I>�n�Ʃ�+[�$�l��ᡣf�����'�v����)"��+�s��!���h�h����Pl-�_�_'�xw�.e�Ъ���Z�@.0�J�Ej�P�vH������]�GyX��0�j��љ���C݂���� �0��ʯ#ޓ���Q=4���"��j��;"O�3�)��o7�^"*���WU�}�R���&�va�u�U�5y��>{C}���]kc%W�4��vڲ�}�&y,H8��
��>j�S�����e"d�Z+�$��w�#x�2�����+[-�,Z �G��uc�8��@փ��������g���N��/f H�OfV�X������`�u��* )�.w=�Z$���bleɼI@�"�hl܅�uR���W:��VzO��X�E{v>l�84$Pk �?���	>��-��#bʗK����O=�%m�K����X_ڻҾ�Eڇ2RPm���W�k-xfyu�%�2������D>�>�Ra
,̀�<Z�<'B�~�`�j��MLw ����Ԕ��z]�,J1ѬI�[�'�1�{��+��^���;���,�s�$�_[�?͠L~���Td�q��lO ߽�1{�:L��g�s��{��V�����%�������2F�f��o���k�\L�%m�9�rA[��D���4�0u`�:���&W������Ўq9��W��8�䇞��l�GC��ܺ�v�����c�\�P�3Y��F�"�L���舍�'�}�|NQ�W��!S����xp�����Zh��c�o�!�r}��zk��eU���Uǉ�>/����oJI?���tß�_7VŸ�'/����מI�V��C���Q.���c8>��Yv�+Eo�	h߅��;ZS,�O��WG�De���g�h"��d�O�z�7��&�x��`���hI:���d�U���e����� ����2��س�M�O��p�o�$��$w���cj��˷���kJ�Q�g�!嶒�@j: ��a�M�f˃������f�����Y�������|������ث#j��F.v����g�هրU���eyL�j�1��ԑ	C��������������{�lPbt;{�b�^��7�<�.M��zV�V� �xC��d3�t�Ȋwi�Y\���b��Ni[4�VL�ʺd�����$��-��j	��f�װYV���uR�������v���y���p�����Gd�'����e��w��5=`�d<;����R��e+��M%��6�Dq<����R!���@����s�E%�EY���*�y�C�+ݡz�|�G��ln�w�!�� Si2�K���4���	���YZ��_�e�E�F�y��'���#���ƪ�q$I5�n��T�`o�+>���ɕ�<ء�o�]�DXf��{���ƱcO��ܓ+}6���Bv aRC�)JJ�����;P:�J11�\�Xr��ݕ=@��5�'�qkW��(+aQG׍��)�>�x�=���,r9�5��*���;���1���Q��^(�5o�,$H�-LjU|�Ў��rA�:ׅ/�Ɏ^����]?�h~o��ke�����F��cݫ��gʥG�6K���7{f�3cI��^�: �F�G�����
�h��+���b����*�b�'|J%L"��d8��=f�	L	�b��4�a����C���al���X��E�K�Z�9�[�!������՞��V6"����m��Od����2�8K��I�OF��7AQzQ�Ny
�T���)H��f+�ؠ5w�#>������љ��y37SPu��nR���I�$�+�@3��!�n*���Ə�?�#j(����H�d��j���gI�^�b���A,���w�aٰ������k��:&%_5�ƨ}v�#�{̪s]3aK-���n���8,�������v�u�s�+��$�������p�g�ִ�j"o܉2�ZY��Ʒ��V����;�R9,ԙ(���|³}��M�B�<��n���4R�X��;���r��"I6rUzb��5G�%.%HTܖ��wަ��z�+q���"�s�})'�Uz��֏�����$�ʛ�6��r9��j�J��K��

J���������c��@�د�H���+�R�3א��]��hy��]�L{O���a��u\�~��|�{�bm��~
�I�)�׏����.Ø��廠{���<$�O՞ d���f|��p��ؕ�A�r�R��P�%� �r���H��M�T���C��//�	�` �s�8��܄v��S�hD����,fߡ�����3���6���$4�t��sٖ�I%s�4iC�����4~����
�������j��%7�"a���X��f&6U,�Ӹ�韹A�3ɛ(�ˡ
�4��dB����U�pM��"���4��]�Le�z5��A-�C�Q(%�<e�&^�"�b�g�����Z��<�4U�ֹY��z٨��{�/�c�?�` ���D�r�2�ix�!�t��{��jX����KJ[w/T�������M��9x-&�4$.a�hWX9� � ���ˣFt���DɅ��uh_�c�|�ϭf��f������.6�>���J��2ɤ�ߖ���I�?T���Lo�d�&]&t$Bи���r�4���He*	�F,o�5��+�m,�O�e�Ľ�@U�m�����?zgB��L�aw)*H����3x�P)8l�䜞��|$r/Ke����ڵR8!�I�AV�y�J'xLY��~!eEM"6ͤ#�h�g
[]���A߯�ڀo
kL���N�0`����6��z�K�r����O]i��e���Ï�(]L�^����7�E�'-��Nb�FV6S����!sI� 1��_���#;NW�K��)֥A�k.�뢿��_�F+k#�f�|��j�ܷ9!���V�E�Q{�������ՓTVU���;6�N�-�[�:�<����ĹE�Y�ygn[SZ+����W�B' �eI1��S�QC�7���GcHJo!�؉,j�e�����N�)J��N�&�������Ȃ\�FױG�A��%�?�C�Ē�{WF�1i�4M��"�4̡c��_�%���`P�[nKFe�a�G�� ~�?: ��!�4a�h)�݊�<r����!�
�_�)!�Edī|,&�����H��n�V�ቿ������}RtI/`c74����Q:q��lH/���QT��q�z� ר
r�6]λ��G��?=��{�鑏����G�~�3��r��Q�y�\�_��=A'�N<���C�������y��Y����or�B��3��:4/�][��H�q�􂑎�L�gӥA����=�)��]g����Z߈�~�����#,����{P=/�_RHE5��l4O�x�+�jM������ֿ' �\O��nK��`i��p���tπd�!�?9�Ov�i��A�������׸7=�A��m���ҥ7F11�=������s�$Bxx:&�_BD��,
3��Z�r���LJ�B����7���5A����]8֮w���Z�_ӈ���!�/֑\�eE	�-
J��ss�B�j������<`ɼ���O��?�M�f�o�:>O4.�L~dL���F���U#b^Hʦ���?���iL9[����M�	���*Uz`�=J�i�n���a�#R�h/}��L)�B��psu�?���>( =������ 2z~�:�ù����C>�[�(c@�9~�,�wwkuv<�%�UQ�G�1��k4%>�D7�4>  b�l�o��V�TX���w@je�7R�4��	���a�EsM��D�neh;Vh]�}��Kީ�aH�Ë�D �<q�'���Al���f?��4C�*/�WV�����|�k�L�����Z���h�*��5L�~k�ݒ&N��. D"3�1��
q;F�X�4.��L8 G�Xfg�R���=Bղ�V��:�9!NlB<D�L1����EW�.�@��fü�S4��f>?�	�O��|��Qz��>}�U�"�n��$R�e�����'�U�xDv����:9���.L�+"�����U%R����G(��;��ᡮ4o<SU���b70>D�^e��+��D6d����Vj�~�ߕv۶^W�2� �ڢ.#:yH��fX�DZ��X�O��q{I��PQg�|O��E6�օ�0��9�h��iv�,�!o S>�R9@d�����c� �mCL����o:�,���~Ok-=��U��ԫn]Tl��7��դ�e�nփa�:7��:1�a��ځ�ӪT�:� ���^���)M⿈�H����x�,���d�0���z�a��S�@JMw2��`85�2�kJ��HZ��Bn{�<�\��*fSU�KQ� Z�`���s4��Ҩ�X`�1��,k���o
C;�1���h�@����⶿����D��p��z�	����U�����q$c���un짜�zDMjS�[D����+��rmT�L������w�}M��~+6���n+:���s����)��RnNe�iB�s�A�a|.-�z�؎��^M˴(I|��]��)�H�w_�}�L�
��s�Wq�I\��MB�$]\a�ƨ|Jtog���41`1T�ƿ_rzhǠ���լ�Nؿ3�U*h�a#�K�W���������8�$��������c7��|��g,��x*B� �)	)���.�u'N��LY6�%�p��3���ǧ{��
;[0��f�(�msq����;`�rN�N�j8h[�y���À��ő�]�Pmg!�5�S�5��7�g�^�[�c�R~fm��������	=��H�"%��q@k!�k�+�m঑o��m%�l<)�">J��Ƒu�e�_�N�%�&[�r@ˊ"����s����w�T��(��������O�Ǽ��;���Z������,�{y���9<���0����q�m��>�CD̫+w�ԉm�Z��T�����,5uzS5�6�e��FҸ�6�C8Y\��ǩ������
����ԿW��AxfKty��݋���i���$��g��;�j���I���!�������hM}V+�>Hjj�t1�:������-�<72+�}���/��2�j�y��!n�&�H�M��H�qam�}���w,9����s;f6f�t�E��>����^�?4��B!V�{�������#�`*	�U��%�|�����aQ���#b1���C�hm$ѯ$�G�)\��r�&%ˏ��8�Z�`c:�I����SpW��
#̦p̪v�O���/��L`�\~�0�|����@Ei�Ja�P��=t��	@�Q������%h����Y�Z% �v�Z�'Z��p�`���n�6ݽ;��yz�0��o9D�6	�g$]�g >j����D��7�1Mbq��m�A�x�j��M�F�S���3��m���2���|�hI�[�����]��n����_v���fj(��'L�v���=2��=�?9�K	*��1�Cw���U�����D(��T��Pu[I� f��CV\ƞ�K��^=m�0���Md�)1�����>�u�R��!@H4�c]눿���c��4�����:��/KQ`��f���i!AՓ�jD�>�@�������h��h��&<Y�Yn�I�_Uc&�HM��iR���ܢ�(��^d�:���M+�ޚ���*=H�R�
o�b���i~v��j�z\�g���R�s_��v
r�����E4����_�c�lh��#���_�]�j�l_7GNuy���E�-�t6MBh~	�pю�����wS*�N"���7K�$�+_�]S.,>^,UF~�����'F�EB��C�N*
 r��8sn�~������ �����Qa�kZg_z�lfܭ*�;�P�l��xGpq$ʤ���@��'�hU6>⤘���c���A�ۍLJ����B(�i�KY.L[�B!x�A�{�;����خ�,C2����RFқR�{�8�K���Z�E�ǀ���ȳ@ �%#-n��Y;r�ʳ=h5$B�M��%���w��ŝm��=bi;�<��c�88��@����C��4>�N�=��<u*"��A>.u�u9�/Lי�(���� �2q�Ʋ��{0��N��_/QH��º�ݏ�7�Q
�����OKt����E����"���ۮ�,�(�F�U٧WI����F��8��8r���V�ڭ2�i�2���|�R Q���V-#,h�T�!�J�d������ J)�P����Q.zX��D���8U�@�#-N�v1�q��b�7͐���:�ue��tV�5�~��=�P�`�wB��� � {=��k?Fr�fݔ@k�r�ws6~j�&��a4��ðˣg��������$�����T���W�QTZTC��6�r*B�8����6�׭�PT�fu�Β$ZwZ��Nm���x�;	E� j���%���DdX� �t��O!��4���J��I���~Q��lOd0ᝎ:n��9�Cv��ĲWZg"������ݼ����tnnC�AO�e�}�{�������*�{�KD�9W��L�.�ܕ=��[o�U�'W��?S��٩�9��c�2��i�ك�.h��ؗ@��꽝.�J>��E�粗��N�}7��kQ3��lwʖ��W!�D�ĽV;�8c���N Y೨HO�m��g������{	Fyx�>�Al�=��b�r7��t�5��q��T{���c�ۜ���q�`�:�I�
�LC���0�*WP���n}њ��{<f��,��9�N� ?�rbΩ�>U=>󷾼�|�p���W���a�l����GV�������V�ڱ"�{�Ơ�^���&Pr�ʽ���r؅>���n��-�k�C
?enC���T8t�+K��ۼ��) ڟ%@9�����^�}TAD���}d����beE��J�oB@bI��?�Ն#>打~(����$%A��y	��
����y����l��<���l&C?���e;�ύ�Yg�������q��s
B��+sc8���I.���S�ZP�n\��6����f�S�P.(�0�4҇$��:�si%��&����A�ޞʘD��K�1V��,�)���,���Kl��%Q��@���MV��}D��!�>XL\7֞K���}|�����J���it���AƯ��5fЄw����<,�r�
��%���Ӧ�f��~5��8������єq!F7U.�Ce]�����r@ϚV����t�Tz�ߖG����t�(����KbX���� W?�[a�X��{�qr@��T_Ë)8A��'� bI��?d9�[8i�\�J�f�1���8�q�e��?Ϛ��Sh���hXS��嘰�����3�4�W�m���^�m]�$���4��.�O�{^i(�S�������'��).adK
2/�d I���Ķ�N�X!�zr��""��EG��)L�G���
"�����"���t��B�s`���$��w�=�+��P@��
W!^ ٙc5�L���W"���T�%�J���5� E.�����ݗ/���k����㭻gߋ�*p}����PaN�;�m2 
o���	���Έm�v�?D����N��e�9SG�q�a�Y�V��>y=�@��r`M� ���t�A�mT' �|�㡗�\lW��%�:�/��\*{�K���n� ;,5ŠU2����9��/��ì�9�0�o[?<�A�$Z	a &dT �