��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_����]ׇ5�F$�,M�6��"�����hgu��:?)�V"*�T��2�6�v8,��Q�3"S�Ƀ���+3ӊ�ɽa�xw�W&���K(�j�G��O���s^"��V�\#ZC�'l�9�C(�N�����5�uߵ�P�=��i*��fG�.�����xvE�Ц�jsLg`.�ߘ��w���Ǖ�z�8q[�Ap�Z�մN�V�.�XV,$�w��8����]ϐ�{��ok9�Ok�g�K��i앿)̢�O"���}]�<�{��)�u	�Ǟ�DE��(`�7���}�[���xW�*���Dh��Vv;9^ӌ���8���Ќ�9���$�*�>_���i|'L�;*=�v��+���e�i�J�K1cO({��w�}�.��f0L����琜m�22xs���5	$�x͸�d�� ���|��M�=���6�h�dq�n
+����w�����?�.�%~�Xb�zW����O��H��TM�����m�� ��Mr2����s���g$�O"'�hy�c�����?�B��������$�w?j�(֠OxQ9�����H_�J[�*:c�;tc���5���s\�Ik��0"�;,
����)��q��>=J0���UA7�hE�<?�m���Hѿ�a��.�A�׺���h�Y1��n�QWb�'rN�u\��U��/�&���r3����p�H~�w��,�P+CJH?��MA����θ�Đ�0���3\ ��k�}3������ʚoc̶bps�h�� �m�X[s�M�Wg��"�y'�@�T��L���5粐�徇l��5/��:^����%��QT�o����K��"8*}�3�|��U�΃�Z4uL����W�$_��m?՚���A�"�V��<�T��+��;��7�JS]~����_�')�~-�ӵ�w���aӬJP������_�5�ny�QTl`�n��1F�͂��
��KypT��֞�#��|�������)�T&#�I�/Ta׎.�̂l�4�0f�;�r7Xf�֔�f�`���P��` 1k�i��C��sj����|׷:�w]3F�*TGr�*U��fL#�޶�嚮"����.�)�
eOP6Eh"͚�z��T�S����HI�y�6-�Vp}�+Q�a��(P{6�La��T*5��������f��O��z���
yʖR�ϟ"ZF���E�0�D���@�J��������ļm��Ӱ]��Y�\��1�}�����u��05�U�! �zҒ�I�r�by<�6^������<Jx�t�`C?��ڡ
P�CIg�Kr���?��α*6ɩ�#&�W M����ۛ�r���W�Yg�	��5�p�u��8@ʌ�H�U�D�}]�5��x���\!2���V�}�b7�]�ڷ,K%��7sb�<O9��1��v�AD6�[^<����4�x��Ǝ���4>�3���Q�+�k��Fj�=<�{E6*�0�E��᪽�pk�` 6����J}��L�g��k���2w�e<��	��Rc,\�� �އ���4�찜%�����6$�u�灾qN092ҭ��=1�V�R���{Nn�+��D��VR��r{�O_�q���)��E����b=�(^G��e9O����;���$~�I����hp�ݟ���fGcW���P�6�y`�d��4"��.���ӝ��W����b�M/jk�� Ux�C伍/%S����th��M� �?�E��(�ϟ�-�~2���nz�izC��L����.�����$+=a��WR���_��h�2L�;*���[�1��"�\�bnt�����?����@�@߮� ��;/���G�xC5a�.�>�lt��*����t72�+��zK��譽���'_$ �:vBB^E���B�V�,�����{�$>_���b�����JJ@� ks���5�CDDQ�h�N���i�
�*B3N�֑pȺ6!ՙ�|P/�^��ELK�%��X��h� �恙�H�m[�x�7�ς��4�P�?H��{\"Z+)��-�ߟ#Z���*<O��_Pq��z��X�'*�QX`�Bѥ�p�#����^bT`u	�1�����lȴ�SeC�s�|��g��M����[IZx(� �lŻ>�$��f莻L��!Ze�P�Ds��0�����?}Ϙ�F�_1ku���j';)e�Y�i6��	��o|�uy��0}"�-KY]�X�p��A~�[�!�V٘�
�)C���?���6^ʞ4������.��\
y�ŷu�4q�S�� �y��U
'aЁ�x9�trnKp5Y�p�D��gqM�gA:�?���4(�S�G��.u�Hh�M�STH�ÍZ��z�NP��~	�����F*��2����hFBRa ��]�l�W�?�@��/>���{�"n�4<R�M�U�zt� _����Қ�����N��Pӄt�4���/pf Q�J�����@����qpW�����;��фL�;-pI�z���Kf�A�;�?�
���wdM+�E
ga��*����.k&p"�]+��z/�ֻ*�S ��֑�K�Cש���U��:h���U?F#��u$�!O�>;&�%1C�߭�RbN��t{*M�
P?Br�d�,��1>�����z_���fI��,��Z��k���QA..⚴�|i�a����w1|n���F#�q�ߗl������c�ÞmI�% @]7�"�˹�u�V(���+��z-~@Z�W��M����>��4W"m@�LhZ��ԫl2
�o�}r���ӂ6����9K���@�����B%3)U{�}׭/�s�1�r���:(r�H��*�Q��ǰ��I�'x�VX�=Bb�3��4y�� �qya�y��
7L����ڰw�8�� \XP1lib���l΁'i��mY{�Z� �b�"���U�|��Q�>1_ܮw}�ߖ>��x V�_V-���.D+q���afG;PŎ�ו
�,��r���Ur��[}�����}F,��i_��_͜���b����M�D.�$�7>��˟$����ٍO^�Q��Ҹ�!u�{�tu0���j\m�����zpUy�6jL�{����^�����H�r�cmK��{5�&P���9�R�Ӫ�b�	�b�����V�E=ԩ�p)�x�6��_ �_�P!yIec��ȃY�b�or������W�1lּ.�P��#x��:�ᕾ/�s�'���|#��dVi��7�V�,<6\���C���H���b����D~:��@�8�JC���y���><�fY�|ik���ow��p����Fr����;G��2b멷�xߩ@��$�˶Q5�jdџ�>����!QF��ѽ=i~�\�x�nZء�����/~���S����ഝ�� =��"~y"�	�Y\Aڰ:%�~cdgf2��1u��i�Q��Z��v�;��Iʨ$ۙvMV���u�BTd�+!ǘ�ۋ�^�cN�F���F�B	�]����,]�Y+����QT��)�+"�E���&��uo�������P�;c�`8��f\Ls��N�@�uH���5�F�Rl.I��
��Π�<i=��a�na�͕M�%,�P��}��۶͞q�G��i<hkK[���<�z@b��7AP�����y��բbWL_��iM�����# ��ؔ��W��O���׿�C�Ys���]��rr���܆OG��h��_��i�����<�<e�p��� l���3,���A�Ֆ6֣?V�y)t�+��vL"n���#!��������kf\z��4,�3��
+uh*)����{f�~�M*Mlx��j��5җ�Ϗ�� ��:��7��O��'�̐�
�6N�u�ܹ�m�MUf?�5��XPR-�<�5�Nů���l�L<���\�7�w���q3����J���������w.V���n)�״�am/�nлA�oo�2��j-�]�x��GB��~��[:��E��i��݊�)��d�cd�f2��CP&le�F9xc3���n��o
�|�9��`퇨��~�=?��
`�⓿�樔��k������g�0`�d�_QM����X?�M$F3$�|� ����tU���}HMi�����]�?���Zɨ���ҲLߨ ���Og����� �i�s==��E��aQ��tn�"9S?�ЍA�b���t��n�e�/^|�,��߃|5(���Է=a��|�?�ds�J��eʨ\n�=ͷ;��ǰ5��Q�&����P@�����������ۿ���Q���B*���ӂ9z�I�ؤ{M1b�ΙO�	*X]���e�j�uIo�s�\B�:��,�n�����R��%�gl�-P�;ťؑ�c��_�`�6�,s�d��W�Nx�8�
#y���KH0��撬�)�/�D�zÚ���t<�,��� ��&o�g6����V�kl�>6���EXoC��2�j�,&W�(Y����s�wx҉�ӪUh������%k$qr�Ub�ۢ���V�����|
s���4K�-Q��"Ǵ�4l֕be��sn�|'���>9�Џu�6����/�%ɐ1 �����V�g�	W0��ڟ�c-��Z#�8�iÊC�:V��Jh=�6�a��X��Dr=۱�h������d{��+h�+���h6��EH�Q�@�^���Rg�K��.e-:.���R�b�$�P ޫ�4;��;�Q[\8.b:�o�3d�ٍ-E����__�9������fv>غ�x�㴈�J>e��G��Qjz?��[t��^'l�;�X12��D\���(P��U��/��w:!�R�\T�t>����V$���+���)-�!�5Rۇ��/��_�M�,S*��(�\��j� ��)�.:6����Cp�~�וfէ� ��<ʚ��Hx��ܜ��0g�Y�og���|-^��5�n0}�����!��P	��zѬ9�����b�K�w*�8%�h��/������ˑ���e*�6V\XT.b{3x�!�,�r*i���F����'�	|@T�*	�I7���"�_W�P+������Q���%���?O�ؖ�(�gq�L�U.�ӟ���{�~=�x	�S��Θ����)���K0X2o��$��􊂗§�HJ��}�+�T�|d��ໝǶ��g�l�@g
��;��^٘�M������7 �ʞJ+���&��(c�,�=�|�Q�ĞI�5#��h���c;~߯���۳���4?%<�v�i�$�Ur�(ƶf����eT�O��O�A���
�Yw��M7an$�>��\�&�4��������3Β8���Rxzw�'K��j��Ak���D���Z�*���~�s:�����%��6rB����4R���f��lA@�j�/��Q A�,P1��������R?*��3��R�� {��	���X����QKk[�����F���}���m�]/_oѾ��ڨgvǢ<@��˘=��J�c�8f$������!�<�����dS�gˊ$�����IL�Xú�Ɲ��%��qs�UD�h��G.ML)���jG$^����ģ�}%\��S2��<�-�ehX��gH
��e�+�I�zp��p�P&�c��T9n.�Y]�`C#(�wNp�R#g��0�9�{�b�p��� c��������\�o�c^.C�M��0F(d��,���rI��N��cŁ[^�Ya��f��4(o�ަ�G�5E��L�)�xV��|R)�,�\�wP�u�_�𒺝?�7U�S}q��`e��4M;KA�{�(�@P�J:M�W��T����Q=;Y���:��6�������z(h���j�s߼�氝���4G���߾/��`>^QR/Գ2^���3�U<a.J;�~-�oLK���T]w��Z�ұ�"��X��$����,=;��PWZyъ�Uc�h��Te*��xG��$�S��(1�	�79OP���P瑼]�?<���9�vg�7��%m^�j�S�3I�6^2!n�B�,WfPߘ<�8��Y%��΋g�9rV���I���H��ZQ �v��k�3�cˉ��X�?�XڭD�?��u�x�:a��?�얡�_r��ʕb>ˣ�8/g��JRE���g:��U�K�`"��Z�o/4��o�ڣ<�ME�mA�qq��'�w������U�^q>1n���9�Ƒ��i��48��_�+�_�{;;�}��AR�@#Զnc�w���t��2�U�.W'�{EA�4�1��a�3�18@��9�Q���?X���f���KE� �a	��zI{�8c	���s���^���BQj;�5�p�ʎ��4�r�ف�����#!�DB�G/�� %���jg�K�u��:��J�Ӯ�ﾦ��v�ؑ@'�)!^3�Rj]=a5P���'�S
���"�=��Z��!�9���!�婺�F'%���%�/��L���Η�L!l�4����X�`L&'���{Sm�<8x��sB$]�uT{��S�4�h����'��뉂�S5SGR���y��^V�=��dT���R.�w;�|`�����>�b��
�x���7�2���&_�v[�v\�� �Q��d��.�.�3�昵���vQ����b���9�ԅAM����+�A�ࣗ ��@l�TUݵ��M��v�_�*�pFEO��ز�������.W�#(��1���S��vk�G���
)ng����B
��{���-*'�?ٞ��9���޴L�7���:?xW�_N�]�@�v�^��Z�ho�M���cٴ��C�D�J��}&�A��;�7^.3��$�2:���!��U5Ϊ�Z���qQ��"s�O5�C���Jd�oF�j�,z���U�k�T������B�0���t-�Ew}ND�	���FU̓=�?�`����qnx���;�>#�7V�X�u�e�m�%�6/�N�ܑ@��1��92���UB��N�9���C���Җ=ϣÌt�$j1��S��Yqpzu�q�)A�%�8��Ū�QMЏZ����m7��N�8.�U]���Ҩ�'z�S!4�N�9��l-���A7�u���5�� �*�P�y��}��|A�d�?��`!c����fJ�Ƹ�����'
��ӳ�[��wjx�s5�j��s iC<JK�-�t5��.1� ��9��w�9�� 4�a�ѿ�ͺL�4��Fn�S�0�3���h�J��'z�(�w�b+3<d��8�ؙ:aU_@(Hd�o�E�ȇ��,H���1�՟)㬔��C��
��M!O�2�[�]� z�5�o����$2u�B�l/�kT2�9��H��;��A��6p)�`S�:"Q����~�wnQ��tv���\}��
�F�a�¬L�2vKw�Aԏ�1a�I7�oa�&(SК^��q��@]O���{� �f$�@���ǯ��� ㊩l��Q8;��GU�~:Q�i%��/s�+K�\��s��tD� ����(Cs�!�z�׵��h�;3�bGV� w��pqD�\)_�T�#&h]㍡	�q�h �<)��'0Q�5��%��R�I�	
4�6�w�%������CD����J�����`r���H=�1YﻇȐ{M�)��^+yo����;0L�)XLǙѝC�,���k�{W��$����'��3r������{�X��6�<��#��(?�ڊC��BR3HC�Eq�9t�� ��Y���q��O٘�]�k�T���1���Pz����N�R!m>�~�aCן����E����PMSu|B�|�C]�d��(y��u�i�\���y��k���o`���Y:�0kO641����<.�R�4q�I��g��@6G��WG����y3�.�SH;�K��˒h�]xQ�b<��t�	�?W
.��ؽ�,�/�kƅ���v)���x��f���MYQ?�6c��	�p�ZݽOZy��I��93��G��=5��36#v�e�W�Y������D[��)��Ŵ<�Bm��|�304���hKp��p`��iP�e�����;K�_��3l�p�
�����W�b�~�S�϶�W ����L���m�{]��|�e��y���Q�5O#�@\4CiT�9H���ͼ�<�j�ߔ�b=���o���°_��Q�V �|I�$��u�вl	� �а�FJB$����A��?�Ĥ���cͮЗ��)�!�K��L���S�!�(4$!o9I��E���'���b�i]m#�'���ub��g̗��c%H˩^�����"�f���b�:6an��"���s�5�bY+���.�3}�x����=1�Y@C.p��ee���G`M;=��1���C�'q����{t���+�c�����'\���揬��C���?;a�H���%L��a�D�~����hh������*��.*Wdk��.$���V�#擐�3?hn\%��O E�y⺍���k_�s�`���5\}�?�C����a!o��^I�k�D�|x�aa����N�up�����^ƸpM�z&M��+Ϸ$�m7�#��:�Y.( ���+�*�����T�0�0����x�e5�l�^Hip(`�*�V�x�{��%��.��R�Q"��&cd��퍽׵���/6�QE��E�E؋+u�Koǵ�rS�.�R���^��j]�"G@-9�ȱKœ�5��|u��LR��+�%�L?���z9��#�Y�]�b�gԑ�1"�t�����9��1!��`�l&���>[I�Ѽ����(�����a�1���R	;/�T�8��~�ә���zQ�Lb�y �v���\z�rB>}7����a� 4d��>Ee�f-�����?�xm?7�7�6�)��~28,��sh�0��Su�M�zp˹r5N��4�'��z%��E4�OQ��ɈGd�m��	szf"q�@D���m��k��
��熬p�ȳ��SB��&ͯ�"��It� Oq���t6�Wg�h�g
Q}Hٸ`ii�DD8F/�j#EU>�ū���������vV�#�ÇH�u�D	���G�f��i �>�;I�F�P��d"������.u�m���b�ǫ�J��1���U(Vi5�?��vN��b���4��>���ôo&o�R�vs�TI�	nA'��I�n���}����������RN�Ɲ�V$��|��f�h���@�B	�����	*����CH=��������J�ĈV���-��	Q�5�3%d��,��G���
�GV�B#��Z�=�mv������W� �A�U}A�-]S ݷv�xqgלQ��_<LԮ���cT�{%lQ�Ku�~ܳ���!T}r�*$���@3��Y~�p��&&����F�p%A5$��.	��%�
�{�#8��V�_D��<���lT�|
]qB�C������w�s$��OD�wp/�1/����N�o!�̿�L���כf�ӯ�]�ۚAz��Z:�A}�d���}XY��*Ai�v5*�_�qn���Jwحx�`p�A��=0xt\�/���,Jc�E��;$\�Zw���䇅��J���L\�X<ʺr�8@�|�V� F�"A�4OlOf�;el5�I]\=��y���v����b��I��|yT
&�1��O���l�_��[�K��9,'u�Q��Ϫ"�8b�`n.�|�}'����Tu)��SL�"��O�32�5�UDy�(�L�Gu��z�������&��w$����J�(�����k�Tb3�k�h�sW�̍=�m��
�g��l���>�D�/�Vk�ҦMy�GY��;��Nh����2=ql���f&���Ad�ax�P�BF6Xt|:c��E1�\1r
l`;`�+C�p�I�������DN7����]ᦼ�;����2��T�����*��\t:�o�Ln���t�_�^ܼ�?�� Z�x����q��=u�����-�7�h7�@+[U� 
�9�Fn���;�l�X��<��>ӑ��(�1hU2��O{ט(��b��g(.�����#�rL�qc{F@�D��]Gsq?�������+q��O��=�]h�����W�q�2B�I�l�4����֙������_�Q1�W��+8���& �z���@Cչd1���a�l�g_?�`�3�/y����~���ޞ٣�-)���/��-�i� �F�L�u���n�����ڞ��þ�7Ģv<-���3���6�԰@X��F�*SE��ʑD_���Ep.~�6N�2Ts|�h$xv���я��h�H�V'��O.��b�2B2sn�8�9�IA�K�d�<OᚧXr��:�&�x8j���V�����8K�Ss\�U5�]�����1�y���i�Oz���R����Qv ߠw-Fmf�Gz��h����[83��1��FbC�wdw��U�ZH1��e�/���菝�5`�Ꭻ}�3�82r������8�$�%a��4R.4�PO��߅���δ��^�DJ������_s\b
�|�]M�D����P��;��b}3��ui��.(�;/BE�0��Zv�����2*�5Ll�0�ReeU�5���3Tݓw�RE�I���|)\��I[�K���ܓ&�� ��p������QՋ�T�}�E3��O�eK�w���h"��u��&���v�u�b�2[�%�����k�QI
^��ڮ!�`M5_zUl��.��r�AX��MB��
*m�6ů�,d����e}�;a��?��,�T���2�Ǹ�C��J�k������ߡys�V]|�'%���lЁfIxh�@�f���}�q��j��!c9�L��]�w2x��Mn��?ףp��v�z
\��?�o�Ϫf�l��w����.lQ'8b��t/7 9�Y>�An�S3��A9xnn��o)�S��Y��%Z��Z �hˇqxf���4��X�+�ܺ�-�y���l�˓�^)l��.
�$��R�2o��yF��%��M�z	�H���N��
��9�y.�F��Y$Yr�c1�Rı�K�8b]���G'�%eo�{�X1�)@W>�e�;^5va�h�j��݋�M�G�d��ܩ����q_'��M-���W�9�W�x����q��{�b 6�N���:���QE��Ko��mJD�䃮0��L�`M A�ߵd�QҦ^槴��Y��ʢ��]w]�v��<@��M\mη#�7W�>�vT7�*�G�:�^A�k��y�d�;Ti����Դ�|-� �HJ�Y,���nМSo_E�d��&5�ɽ.��C�˻�:E>J쯳���p�n��QfA��	���R�!���N=��b+џ !�&(0� )����x+gU���|{<�Ӟ����	�U��Ҙ�O��t~Qv���ob�Ԅ��J_w%F+�%�$�
�p�9a�`g�D�R�X�g
��*V/���L�O+�M���o.��{��3�=ξf����_����5\��7^��݃����-C�(�� �}�/�W�a���/�,!�PQ�]I��+��;�N������Z����N�>���RZ�f!�JSee����_`�I^t�9�w��#�f����愅�C��Dm��-Z�y8Ƥ,��I�Pý�j��Sث*��Jf|�&$b� �[��ä:��e��_�>�}N�3���O�Su̻����8�3z��}��@�Fk\q9(��?5�M;�������Ot|�Ѩ���Yhʼ�4G\��Gn���CT�%ɿΟ����V^��r��UP�Z9|f���o-��+��C7�'�(�Gb��5�ڳ	ߘ�C�q ���ڑM#,���f���R�I�0�F,�o"n�)D�zD�x4n�l U��������c�I�PP5�	��k�Ȭ"��Id|�Թ���,�J�Ik�L��Ư�H���&q\k�:���QhFއԧrq:�;|E[�B&�"fg�i�~S�5�r�6OޣR�t��A~PZ��l	��UUi��1S��bpƙ#x���}��ZG����B���*.\^S�]�+��ȗ�V���'z�>��za$�c�
�ܺ�5�M^f�#Ҥ6Z$�ta��L�<�|�M^���7�����/P�Ϟ�wb�t`�V�L�x!�Ugզ���7C�Q1�~�ַM��\�͖W<��·��B���-�#�����in���m�W7D��*��WSC9�BZ������6�Y�?Gen� `ؘ���)�%�m��C�S���5aK~\�5ֵ1�� �,�ϲ��}���� �[e��~�L][��nt��:�I�̖dݕ	�/�mˌ�n�@+s9|Jriů�l�} s��ќ�V�;{j|g�7kdH���?,
����ł}���4AK�=v���{i��d��uݝ���V�����d�p�م��;��tt��(>+�\KIH���p'9��i�ȏIu��i@Y��ڌ�����R��NI��.I�ɥ�.b�Z�1��z�)-�����q��@{z,"~�X�����dʉ@S"I��7F��cK�t<H��~����+G���h�7��vOڵ�^B��1(|K����:u��»~7������L��h�����k���)�K��6��ut�7��`��A�a�R]�:�ձn��|uP,V��AT�Tk *���p���cz���H0E&�O����wo�)#Ё��:�c��Hr+&Z[�k�\&�b�Ġ�v�I/V��f�j;����5�7t�T���E������B��V��Ҭ=���r�r61�o~�;5F%���~�|����"M����1���s���el5����5X�w�Q��{|AD}�ȋ#�a�\���dK�s�(bX	��>�û{���ʃ��L�6�:��*y�!�������mN�%�Ǣ��C���
-o�v�x�����[�ЅR�0��9?�N>E}@��
�u��Z&����C��~C".���zL 9m.�����94��Cݡ&��q�l[T���Q��оݯb`�Q�Y���M3	C˱-fj�I��(����ٶ�0�f�h���"�u^�G���z�-��zp��c{����!��u�m�q+<z����W����⤼�x^���1_�S�x�i���eLVh�kN@�_�����4Ubo�2���<��VgMIKD�1�Y�{o��\^t������rg��Wx5C��l��\׽��� .~i�R'[n�	TKB+��ͤ ���QtM�i�}Z������x�.2�a�Sw<y��P���n xe{�L���NIsNlN1+&���퇢�Mv8��"QI�[%��!����w;��SU����tc�^�h���i<��ځ:���0���V�)�r1�V�7����K@݆yڡ�#��-7�w*�%G5m�06Ɵ!��s�H��W  ��Ng��q�y�i�bA�GW�"��u	��_F?�1b(�N[ih��}��ѭ�{�a�^�_C�\��r0�/}~�
C��T�Ǿ�cE���œL��>��4U�����L�	�T�2�ĻdO9Y�ǜ	���~)�ny���?T�[&-.�9�Ј�'�4����VVo�u��o�ز��p����{N=!AZ^������j�@�E`��M5D�������rj��]Us-;e����_]�˸h��<p�n���s��/n�ſy�}a�&�s[����̋t�t�����U�	��sӇ�*,�͙,��i~�C�X:�j��ז��R��5�E��+6��`��E/r-e�!�^yƇW����R8�qmDabڵ�~T{z�t��H�m�f�0(ְ�݈�=3����ݡ������2��dJ% [d��KA����2�6尰D���-�|���g�.0���?�����KĴ�C��Y���G�5�S�	HS��0Z^]�iTX��;rf��� ɶ�*H��j�u�b���ّ���(��$)��bˆ��WIM;9��Yӵ���z��/��V��'����*ی�	uj`:T{Q���0�}�?O�Y�;���b�xwP�y��K�w,N���(
4�-/M"�e�3�d�4>�!���()����]H�{��{��R܏�)	�����MK?�]��ߓ�E!!�}��XЮ,���_�Q����B5�S6����]��.:l�H�d,7Z��(�9��P3�
�Ƽ#w���c�<������W#�G�O	���ٿ��<�S�q'Z$}�.�i����x]�%+*Nk�	;'}Y9���D�42U��}0�g�ޱ$�_yC�o�s� �����>f�n����M/�8'�o��-�lB�6ٞ�@�Vf��
7noI;�\ }-L����o	�qϿ�FP[���x��R3?�X�jX�c� ^��3*�Q�gE{��?���g7����tJ�׬$����^���3�<��F�W�ԗ`��"Y4J|�
j��!�D��ȇ�����i����p�u�!�`r(	 ��o
������S}I{q�A�b?�	}о�VzB�a ��ƇJt~��V��lk�%�;�1E���oEp�1}�
S%y��ܰz6�XTH�ٴ\D<HK�+�VL�����t�a�a�]���i#���N�-_v.��N�� �b-3U_�G5��0��G��SJ.�|�{����\rpx+�ک��{{�4;��fIs����iT�:𚔘�y=$��ptM�˙|"-�OWW$R(B��V5�8I'_3�P	��E�����+T��\,�]���^IWͱ���s�R��t��`"�秸Δ~"d���T��go��'�$�_���e{8�L�3��l�5 ޭ�K�Jj��͊�c�>w�&����;�F �>����'ǘF�b��υ��]�_.W�V�.��ݬ@�j;}���s?�E���eM
�~��[Yz5�p�~Q4u�Rdb���ϨGQ���V���c@�}���#�FZ*A�n�X9�W{��My�;"��[��ً&�Ǳ+�����./�Uo��J5W¨��^/ǲ�H��N�*y�;����\�ai�h 	n�V���!��jQ3���G���9/�[�1XQ�sh���ݫA�� �5eٔ����Wԅ^B/����Q��D'|2�s� �۸�=�,�T�т�I�7��ﭙ�r��|�c�J�C�h�J���L�v+���Vj$����mY�ѼwE���ܒ)�#�;
��	.K �$o�{�U�6˔��>�t�P���Bg&�&�K������oU���$�]+�O"���=��ߢQ��n3#U�6���,@�(�1��m|3�
��י�GX��j�uN~u�]C�mӘ�� �*�K��A"##�����H��r��8d�I^��H��2K�o�lP`^�b�|>��B"�
�y�g���.��S�#���w��#�������Y.6��SN�x$��}`oR��J����4&�_�J�P@.{� ���^r�J���<N�^�u'�k
�H��w&�1��cV1Do���̲Vߗ�Q1{�=�͊��:8~��A��-����C�|���fʦ��q!��L�znV��ֺ]��I��r��J=i,�" �VG_b B�Z��M{��)ļ��A�����F&�%H����m���^��S���Q���d :�àɴ�0ǂ^���k��M9M���TG����S\>E�n��w,��\��1�):jc��l��g�c����9�8�+c�,�b����1%�5s(�%����|�!"����SZ����Xw�C˗F�S�d�k-�@͌��_��w�Psc?_[w�q4E�6Q��N6n�۾&���|ld��>~�I�~�zn-�� fhf�;ya�A�]t����A/�'&.�Q0���j�
��?��/���7���b"덙1���ʞ@�]#�đE��X �z �
�!���������j�G�N���x\u�sVf�����;I8�h����6և��r[S�9�l;yԪb�C���o�&�Z������1���ߏ>Ia�y��~����-Cm��&�t��D��#�y�Þ�3������� X�2�	 �9]��n��1@�?���'ޝ�{������W��*���«z�k����mXi�jfM~�˝4��i���/E�B��X�Oh���yԅ��G����������[�'��7+*�
�B����|�0LCϭ�~~��w�0LM2�T[��dWp�&
��@#l���"����1�>�,ޠ���#!��~֝��^)GΩя���
]��\��_��_�F�����5,�eA�I�� ��P�R����gq �P���6r��wg���S���~�$;b�D�9"2�oռ��,M*g��|��?���<Xɍ���JdQ�+,�EG�6 W7r�eyL�?ޣ?he\��֐9M�t�mM�����F\��/�kR��!�Ϸ���u�:�C�5�k�AgR�c��-��iz�8|;q��\���%=�d�o��~���WmH��
j����x��l���� �cN>�������	9�PN��H�.���\:��[�z�-h�r�
�7Bh *m�Y�T��}� ������X �%*F���9�]_s�\�Ԡ9��/���9�M��|��.���z�a������dA��/�*��X�F�UB��Jn�,Pҡ�jNP!����ψ&��Cw��&?����X�N�g:����S{t���[$�N�E�'�;��O� ��7�+�}��\�9 �ш�ԣ�K_Ҫ��ԭ�0$O.���u�庖�j������Z��^�V ���r�q9������3��Ʃ.��iy��� ��(��\�(#̘��^�Xc�#�ai�=�`n'�b�\i�!n�=��gH	8x#��.S<�GҒ�«D��^d��mw��J�:�q �}�6I8�DH���2��5��A6 J�dX?���I@�DH�e�лZ�^��@\y��F��Y^d�(q�/�w��uz�Xo@
>�M��S��]�p��+�/UsD�䦛�����`�^��s!�W�sAS�����d�3'�֜�D�*τ��3���[c�G*�ֻ\;^�Wt�ߤ_4�����j������L�="6���U�FLbm��Ȭ�5���C�M@�Pc>^]�Q�� Ǹ}SYs_o�B�-g=��)��Pn"̤?a���-���\}�Wy-t�Tĝ�5j!��Rh1U�K ���hӫ�<��Ec��
���pӛ�e�&��[� �%���&�_�v7����'�CA�V���\��*S�V9�{�2���P��?�d5+��E3���5��^�":kϟ���k9(D<XȄ�lp�N$.����Q��@Q5�Nj=�'T`�������^#t���d��4�xCf�
>��:��b��˔VXq��a�����m�[Mo���8Y$l�A%IO���={���Fnx��+���~��38�"�"ФZ6���J���jf��M�[��7����jz�m��m^�;fcu�_ O��z:໘�àNU��"��i�M
�S�	��y�o�g�:C��W�8>�.��� Lxѕc�w��m�x�+�����ۆ�à���������;�-�@��2�Ë9�F�'~��x�Y�g�J�3R]rR͕�R��rϣ����-���,bm�bK����Ƴxɇ�������Jk�myUxf�)����N�d���-��Y|P�b��S*��ǆf�1hv�CA�������o��vtJ����1�K֎����Q�|��v�*fB���;���\��釛���k�)[��^�Ӿb��1��ln�	t3W͜�^�'��[1Z!��jBм���Nۉ��.�vV� &��Q��S��/�t���*+�r`֑t�^Fx;u����2<<��)Fڱjɿ	[��\�H1L�}r���<�ْ���Xu�~�>b�BA��
�$�8j�eҵ�苢2k���K�5ŗ��i�}����5�[#�kp��G��1P)�������t�CXp4�8	�B4�%O)�uZ ���A���ZL1�PrB���a�ՠ�5?�/?��\�Jl��uS`vnmp����J���f�j���9�-�8�nC�s�%|������Yߵ�fE���W:�����W�?�$��!��u�_(+f�ݡQ�������'�U��z�?QY'� ��l�9$�P��"�xKH�Ɇ�h�AJ'����U�^�4�A�B�Oc\��R1ht4��<ȗՂ�ߜS��,ȉd���Ot��~;n��ɒ�v*r�M=�>MUQ�~-���ҍ���)O�J	G�D��pJ�/��qy3�l� r|��4�
*m�n�W��I�wSޞq�0/���t;�Qr�yC��D��>57����z�*@Y�݈6]���V��Z�Iՙ!X<pXr�]`��%�B0�֍L����z�Y�- 0��Z��8y�	���w��8�ϗzٕ�d��͔�P�sO�<�u��=*���*�gܢI ��~��F�z�◓��ˏ��9mO��S�J��/�̆�T�����d�&i�	N�Z'�y���n�&�{�(~$jG����:��4��ژ���-��t����E��ow���DZ�}&(;��>0�.����M�?Y5D��m�=<I�%:��,�b�Q��pI����U9�M}��������m�jjY
vv$��L �ޝՔ) ��b��|�Y�6�I/�$^���	���bj2!�Ǽ�R+�3�]ŀ�Ѓ!�jMH�pe�dF����j;I�,��	ș���A7L�^��L2}+Y����bOqGf���4���I��;��Kܿt���3���R��
=c�%��o&�ݖ�$��~:�_P@�W�E�W��*^N�BQ��27}��B����-����P>�U�_����X�`|g��<�&�'
#� ��f�	����!�a#�J�L�xL��6�O�"p�'�^�53�2C�(G]��!������u
�7"S�{`wY�V�!�N�Ȩ*�2y/��0��&��6�:�N'j�V��	}�s�����3���������*fA_ޞ�����Hh�[�;��/ɨ2�4���v<2u�q:��s��߽�1�x�-Ϣ�#�Gh�kcV�'{3����8lG_�
�n����T,�
҂��q�8Ĉ],�aj9�Ek�i{���R��y���hH ���M�b�*��<�h���gJZ�)�������l��u/Cfa�m՜�o{�hn]�a�L��j���9"(��(��	J�t��f	�/��j����;Ҽ\zF^b��Y��3���P�wK�y���5&����m1�w�%�4��[Gĭv�&�ɤ�a-PNZ���E��U�mBv5��4�]�p��he
��jé���#i���v=����ө�о�3�K,��8�����u>�߅*���TB��Σ=�[(fn��~���E<�d�Gk�Fg�KV����"B� wH��f8���5Wf�������ζ6�'����<Fq���j�Bk�#�S�F!2��I�j�Tk��q�H��Χ�T�!$�'jR%i ����&1Od��F�M���j�R�C��hs�!���?�'^�P�ʁ'�vR�c�ᙟ������2w�[�?C���Y����c�d���j1HtC�����/(֙���Ȧ�@Qzo����q�#�XC��B��yY$�O&�[Z�x\!�ش��:�����h���\(�p/��V�w?C�D��mr6q<I^b:��v�=�}�=Ko10V�n��΃�s��Rv'��{�����g:�)��\�h9=3�X~���94������C,�݀/�?u�o��db�#�����<ea9���hl6P�:6���x|��¥zv+�V�9�䀲F�HKܤ)��Cn�H�l�7�����;�b!�q~;��M����<�,�%�G��0#��I��Č�8��Ѭ;Q�K��,IP8$�2�~rʙ�p�
�\]�P����@V e]���`䝩tIC{� E���/W���i�	��A`}"�o���r]�w-Z-��C�xM�q��p�����:����ez�,���<t��D|W�w׃����=������qc��Ǻq ��0U�=�v�X* �a��_h-S�U���# �|,P�"�-ܼ����K �!*�/�/,b��^�h2!��e�#��q�>�.C�Y!?�S�Ms:2|�I�%���M*�-���[�]��=�7�S�� ��!`�=>y�d�@0f��i��@����ux��������֯� '���M��v��J��b�`��}�<����������z�b-����b���`rx�9z�~M�i@s��+�H��d��O	l����߿n��f�O;�f9��?W�ވ�>%y+����N���N��6.���P!gVa���h�g��U�Dv�3��D#F��vf��P�����NP���(v1gE0�$���,^�yT٬x0�-3�R��ߛv?m[�zȟ&�AK�.<�P���{�i�3+zk��X�����~5����W�]��3����f/�V�F����K?՜�W�	>ʃg�j�*E&��P�$.��I��4G�{���9*u7�Bל����~
���`aT68����<����ꟺ��S�s;E["�⨬#�X��4S@ ����\xj�sE֕%]	���2{M��L���B��m,P�	Xc���1��4�S!�
tf���P�h����sذ99/�. 45'�qo�����N�}_~��D�A#�&\Y�aӗ�;��MYXBF��o����U�>31��0#�.��G�ec$�Uҷ��Y�S�J��b�|�Ų�W�,}J@�a�\C��a�,�*2i���!�"�>�?�K����}FѦE�ߗ��O/���d�=�m$w���
hf�6��E��N�U�����6Ϥ����9�|��Fo�m��;��a`L232e��<�È�<T�t!�2JT���w��]hUz��&@�qmK�ʟ��X2^��ɼ[����^���u$)U[b��xF�	��tn��X���`�6���A��[MG��Ӏ9b��%%H����X\��f�]Zq�ԱX��;�Ũ�3�Y�nF��%�H�_}!2}Jڤ�.ĐA�������B�T*��+�ă�'*��:7HNW�SU�ߵM� �
_���G�Wf�������8�F�C��(�d�pIv��=��X`����jT�y>��
$�V*���j����*=��'c�e��M_0�� �A"��n{ ��J�z��Y�fgü�Zi�$�N��������.�Y�1��]nx�U� 9�T��
c�d��g�.��% B���[o�C�@,C�ꄜ۰)�?�bv�\-}�g�8n�H�*��0��1��4��8:o��1�ɳ"��bFܛq0`C}s��f��������T'iL�F�c�ȕ��U�nW�b�����󙉳�5X�'��wa+1�����t9\!�LA��8֪���PV=O�d�,c�f~=�+�?˺���:=����K�8�-��pi`Ź󹇟�|߭&�`��c� <���
b�ZJ�W<��f�rm��z�9�z��4�_��4����C�.C��F��\!�����V ������|ߓ����R�4��t��gcj��ہll�*U��L
z�/!>TR�9�I���gd�W����2�֡��"���o�P�mҗ?>�3KQ��x`�ȇ�x��;IEb��J����'9�>͒�vT��o�M��0�\ʀ,6?��h�ї���R&�1���Q*?�����n�a��X����ɉ��#rVc+L겺�� ��e�A���-��ώ��	z�~�Ե��̅:��T�����!R;/��2F��@�''#�qu�b��Г�Q�����x�k?HB��EF��X۞�8��Tp��ep��)3K*Db�p��㴪Ѽ�����@����%��,Q ^����؁��Q�y�����Ϲ��[]���Ǳ�N�W_ԫ�Ll�&�b�~�H"z�m�I�J����(��"ʗ[���'5��V|�6��f4�2 gxT^�.�U=#���9~�3�y�W�Y���lɇ� ��`�i�G�x��������:��G9��0=��v�hL�������x��͓�;�lt��LsȻ�wլ3ԅ����4:#�:�BD�b���o读��J�6�v4���4���@��������������MK_J���!�#n�O��qf	�	9��np�T`,]�PTn�Xյ��ǧV(��w��e��B�  z���v: ���kI?���1���F�VGU��H��w�y"����zpR��do�lp�*�ΰ��s'�;Ly�M���$����!}��Q�9Ɛ�מvM�|_���S�qu��	t!j
�U���3�����az�>5x4W�m@�3U�6��I��� @6�}@,Ç>8"Q��)��Y��2r�O��}?�p�K�~���A#���[&9o�D�܂�m�7����%#��1Co�j�0(q��#f�-�Q�%U�&ʵ�4�����Y����Ba&��������-�[�Gp����a��"��%�zXo[tD�t ,4��9�V#�E`��$�rVFm�#�P�� ����V(-�Ys�Iʅ�8h��ck�4S�Y�n���?\�W�y R�hNE�p��gBeQ�4A����Btp�8T��Bd ֵ����/3͘w�,Xl*9^�&�a`ZA��4-��v7s���_)]��H��EW�0������K��(�uݵ�{�oo8L�=FVM$�[�m�۷2��qh���r�����)5r�m$�َ��a�VQ8�{������,>i)kD k�I-m����we�کk.�b������g��8KJ����}^Y%J\a[}IuB3��cm�$Z=W�������ǜ�ib�T�N򘉭9;����.Ⓖh�2~��������B���=�i�Vf�_E�'���+�7�%���4O���6���2^oi�uN�,oZ.4Ҁ�%s�ғ0Z	U�Gvy���ϱ��<�5���p�;Z�X�-'[�zX8Ҁ����1+�V�s�)��я�d����=��m��=�_� KZ5#�|d`�T,'_��^�Z	�P�q*����Xc�jP��u��d������F��;��C����I'���y]����2if�+L<�B�a�5�`!V�1��T��4U8W�d>�#If"��;��ꦴ�,q���D�5�^|51��	_�F|u�v��In����&��w�{!~5��`q�м��Rk���d���8�9����'�@�3C����:S�)������(�\��5nQ ���66�����Pr�d����p�����*<8�r'��G��I�`�+tւ�Ô6�O��$Rg�[�NٱW�M��pS��[�W��h����h�X��YiG�k)�D9��f�s6��RL���.<10y9on��"�QISFOÜ�:��`�OnOo�K�C�?&\V��� �Xý��Ww��ǲ�ҷMoM9fqZ7Fr��6���)���=D ZNX�4%��R�9ܨU�Ƿ��X�Y�����o���������rj���]��v�����w����I� w����.����^�`x�?'�=(�ju���%�Z���:�W��>�|�Q��ԥ�@u�ώz+��+��*g"���q�:gu��A�ḬQwb%o򻨥���Z���(,|���l�ɥ��Bq��H9�!&Yz� S���c	i���)C�o�i;ҁf�7)Q2�W�� ����\�
�J/}�)⟞��.Z)����y��_\x��T�wh��cb�␞�����
��Qy(�#�$�6�;1�L�����
O�лsFȺ,�0j����ۤ��mn+��&Z�"w/'�&�>t뫴]H�V�v��ea݄��G[�vF�%�F�W�_�	�^��2���Z�/īK�/
)�g�oZ�"���{�\ lŇ�#��ʦ�B��?�޷�R�t`��)�ڡ�p2��T���3G^"Wi�OZHl	Z{.x����jᩪ0��~D�EYcG�}Z9	X��E�7�S<�������0��s����>���*y��;�m�o�N�+����)��`k�߄Vډ>
���r4s��x���k�qy��h�1�huh`�)���V2t�����9'LR��s&��=���-��Nc�w���Eq�v��>�/w�5�Pކ{���*ȷ��V��JT8^���O�orr��O�ӕŸhg���6y��x�4�1��̫14e�	��������i���sj�fNC7�uͫPB��D�U�D�l�����C�1&e�+�{ذ쟊9Zǌ�c1�z��o�ԥ��0��H�4�[����'���MA&j�J�o��ķc��uţ�Zџ}G���<��l�$KD��y�yϭ���^�aN��K����m	���E���2�`�������<^�����KS�:����
`vd���(pJ%A�:����4���<��h�B�c<�`Ɲ,�s)��$�˼�y�O�h�D��);�4���5����$��-:)�f��V5�3)�`Eu���!��ct�M���$���O�����v��C��B��m�kB+��*|�O����������±m�Q����G��4�ԅ��J�~�y����b�=7���ʲ�^�S�O{��G��
������Uv˷�˘�w�/Fg��qϣ���97h�f�ӄ�(�[P��瀈�Ⱦ�����v��W<4�jhpaY�{E_^	��W`�õ���e`���P�,�,��ʗ;&���\��7��6N�ld�qZ����9�Tn��p���cO�1�1R�c^	>Z㹲�6Gb��b�6v����Y�joj������WC�S=��Q��3-��vl�0�\9)ibA�]#������O0aV��*��ܑ6�@�cI�?�Xs���D���g��j(e�4JOK�'��X�ӫ�0է
��.��w:�H�F0��͛*�������*��+�n�`� Y�SH��a[�����P������f={�t�^J��hB}�2�j~��ʍ�pO�1�"�i8t�;?(zw"����ũ� T:��i-��8ʞ�u�\	����R��<�-.^z��e����ktcx���x�(CS[���gY�T��,�K�aH�t���"kW�F�nr�ks� /lt��iAR/�L��o5�35��ʜ1_�]���v��d�tN0��XК��A�eSa�1b��'R��P���B�E֘L��)2@9�@=Z���;�`о�6�p'� J;�5��ڎ[�s�^)䖇�o���ң�z��s�Sz�q��5��ć-�e��x��M=�e���̈́gT�!�T�G]9�̥�o�?�ꅸ(bH�O��V���x�-fc��C�%����1|���n�T�8�	 Lׇ�j�ɓ�,v' wQ�(|�?w�3A��(X���Q�Ka�v����[��Ӈ]5����|�#�>�����UMW��#��)�}${z��=,����}nw���nA�G��WO8J�}91�N��=�F��i��.��g�`6�Om]�w�w�����!�疮mL�+���-^�`2'��:��Q`o_H_�K�`h�t�'�	�/k&���f�џB\��߉��P�I�"�A�M�ϼ4���㍯J���^va�zo+� G�uh'���	�DȾ=�$X}�CD�������[�tL ;��
G���?��9��� �0d5�}�sRn��	_�G�[�w�)��6_U����$�fE��<�]ا��ml��-��#/����6ƶ�K��Rt/�`�JC���RC!��i�	�}�Ԋ�_)��bMy���V�3�7��䱁��J�e�%��`w3���m|>v��!�-_.<�\��m(A`BY���W�#�n=�-��c���������r#ȭ/m��Ur�dDLjD��G� tx�KA�R	G��~��6-�$v��>�t�/r�m�XҒN�פ4K�4߹�hɜsL�����cV:u��b������ۤS �d������B�@Q6i�+���{�FP�|��f����ݡ��-��U����m������T"Z� �0���i�!���HL�6z��Qf��,詀��]Z�:9�rI;�*-o����{�PpO=��ƌ�c�2[@�Tok������I�v�&�L2�����KS�=VO�$��(�s�v*~����_ ����,5��l���`����A���+�K�&�('/�+5����ղ�qے`��_�[��O�B=�cn�~wh�9-��s�;��+u.O_�a��ڢ�A>XR`��������n�#��H�?+�%<��҃�^E�c-ZC�5Qx�9b7D�ј!T��-}5�7:˙�7��`;�D�̟a_|�u2"�Wg��d+�����ژbl�.��j��%�vQ9f���;�s�$�����q
UCS)9��.!.ry���C	t��56�,�U�ɲ>X�����^�e�9f[٧�o^cW��Q��қIV���yӠ��g*����2[q�g�io�3�&,*1�_e@�/��̀=V�{&K��;r����p�2�ac�i� ��<)��!����{�~tp����ު�-ą!����/m���f�Ωԉ.i-���D�� l��XN?I�<�4��h��AGqiB��R�
�|p_��V7.�����og6��W�.��u�����Z�1��Ylq8�#��t��=F�L2���B�Bv�2/,:K�Ԓ��(�9�y�c��#pπ������A�fB����ї�)�~M[+�2��.��"������㻐��� ���Qz�,k���~.���l���jj�Cʰ���k3�K�AS�
.dU����_C_�-{b:��h�O�(��g�`�8�@n��R��x��ʜ���n�q����Je��v�(���v�(0%�����JVq���� �-��A�꜋�Z��3�^«��A��4�0�J�p���C��B��<2�2lIyZ�Ȭ~�q���]b���͍����';}F&*�U�����(<`X�Iv-���+}�}�i6�X�YX2*���<�����Mw4\�fk�ڎ��i���X<u�yl��#���/�Ϩ�
ƀd.�64�>��g�Ou�
Z�Kٝ���X'd;;��Ј���=�q�F��t�ͻ����˿aK^���4�P�+rm+��3� \C^�	���.�V�,<E��[8i��A�1�/����V������=P)�sԞ��^����=+F��S�G$B���c_"�\a)�uW���-�M�� $��U�	<6�7���w�7�)�$~(i�AW���M�>��9�0A�)Z��kʾ��ĞV�)3g���sG���Lr��ӽ��*b��_�Yg���٨�ϡ��,���XH
��oR�)pzP�3�H���s#�yJ��&J�m�+n)��B0�Oȫ-�l�
��A��E"��W�|��jCX;ܪ�����Y\i���ҩ��󄦁p2�0g�T���7;5}�,���Df%�i[mv�3+,�N�l%v\�hec�E�bQF�qF�n�;�Uȕ�E�����P#*w�mZ�L�t�~W�8v��|�f3LG7j�aǢg�������!m���K����<��@�I���>�3�5GoKGm?�e��`��q=F���|��0e����:6<p�ȥ��1�/hN��N%*h|;�		?�ʸ�T0�o�рըQ`�#v���Vˬ�5q��|J} ��bM��>|ĕi�����	V��`F#�6;�_DǙ�jW�zu���&���x��ra���R�ʨ���pz�|b>�NQE3n�{kY���o�"�9t�6�P���x��Q���hG^9�-�]��P3�m� טm^�O? `�a�E!�]M�+��Y��%�׵�/R� D/��~
�i�X�-��Xvަ���[8|�_����q�7oM�^�Р�����~7,<���
����G���YL����)Ƈ���Z�O TV)��
�7�vu?��L"��>��ڲ5W0����a�r[ӛ�A�y9�(W�o��E�u�+RD*'�:L��{fZ�����"bl?����FZ�bq�;�ɗ�կ�Lo��v}֠���t@:�sF 7N���+_=��2�e_��_��5��|�V v�@#�=X�b��'��]/��6[�:t'	�K84?��-fB�	z�̂�� Cd��6�<��*f����]Н���Ճ��%Evw��\WH�D�d�2��ͺ9j�]�\֨��mzS��W>U�i���N�j���\�؋[�ʕ:��t�]Kd���x��{��>^�S�0������3��e��̚����c	���z��,����8?Eֻ��&�����,o�]Ȳ�ꨉ�%1C�����&�#C]4��(�~�=v�6sw��/�S#�*�_��16tY�x��G\��˯�`Ns�t��C �c�u��d�lC�l\�e�崽��U��G,`ΑTk�.��I#6V�)5�Y����#�M?��,lZ	z� ���-*8m" ��A��&)Kd5���e]r͊��Ǐ���'e:~�.k�~R߶�A�\� I�t\���c�LR���q܇0C;�> ��^߂KؤBȡB����o��57���r�LN��X���(\W�N ��}6IbPي�˱M���V7�pz)@ $Z^���u�S�����9-���O���/�`��lw��DGpcz�z��5��o��2�K���u� &�L�>�:���h!o��*؝4��jn6h����3$�vObd�[)�ӹ5*Gכ�����4��u��10E�	�¬�Gp:�Tp�h��`5���en�U��m\�3y��O�Qߠ憘 �?[�^�l�2ma��̭1UH�F�)��''~�#��LҀQ��;#؇)K��aԢ��6����^�B��h�A�a���Ԅ��+����R5t���
0eQ��5_1�z�YE��>���[��S5g�T%a:�|t����)+�":C۔=-	ϐ�^ɐldʼ��hln^� ���Q7��i��?F9>~�̇�9c�1�K
����n$yr$�YA�ܞ��*�24x*:]�&²�+��ǫ�,U�Aa��c=���M@7��_Zc�!i��a�3��_��Q��k㑕7�S9�E��W�����}�M�?m�B�s*Ԙ:c�o+U�Wt5K�*h{��W��b����G�?�ؕ 5ƹT���c�4.�t�1P��V��Zo'm���]0y�1/����i	o�x	d�f�l/�8�oIj��>Vn���,�0�q�y�Yq�3���6���"<�ZҤ�)(S�Õ��U�&�zx`�e���P{�5�Y�D�}o���c�.�GJ�4Tv���{zÄG�w��0��H�VQY��+���C�g��~��{�-
5�M,��TU
��H-J�� �P�� ��M��&��5c��ǁ��6־I��EYULa���+�
l�GЍ��Bʑ�pG�bf���~�N��ֹZ�K���1>ElC֟}O��Z5~�e��+
����%v�R1�����囌&������{%�(��/%tfi!iz��j��6�sv� H�s���D^�T�����թ��
��I�ST�#�����ːN&�6�5�6Pӌ���GUUH�`���,`GAc����}��8���ך�� �"R�V *6&�~x;%RR;%%�E�Κ�+.�^�����t&c-�L�xG��z5�ZؒTz�"(����	��Wp���ó[[,1�]��03�����҄j:�ٱ`���4���:��~�<�D���'^zq)�����Y@l	��Yp����w/�$�����ڌ�J��]AR�F~���	�l�h���}��Ew+/�0�5����V̪b	�N
�h��s�-�\��J��(�}%{�����U 1��<�N%�a���U
/�w�%O0+ݽR�S��7�ɽ�Hظ9u!�w<7������u]���I�Z�@Q�
]� O������#���k+%�t��rw��1��ȧom�Ҿ
�#Jd���'5�>�w�A���o�lvM�N,�i�YR��w�oY8��%_�z�gW��A �^�՚�Cc����W�e(�
x-��	51�GVz7o8=���5�g��U�J`犌��l]%���E�48�1��F״ͫ]�Q��6�����'��?��K�O�?����(t)O��i�叓�aXH��b�=F���Vω�}������5e2���u�\\`6�V*]q8�S�ӵ�$��I�����ALJ�x㐻(����ǐj�dNq�����Tn��\��V}�2�S���D��5��۬�����b8c�0�*��V��[�PW�'[��D��k�����-t(�UY�ƞ�!� ������dlh-�˸������g��V�H5�>~3��E#������B�:���r�1/������l5����C�u6n9��Pװ���7�$��'�)��_�:�2��!�����|@�!�Kw����I���U[�n� ���dm ���L�'��U(ӟ�6���6���1�yml�K�j�1g�〇l�9?��
�Sf8=m�w�ykl@久�RV �F��C����z���RYA��+M�c�栞�R�>�Щv����?��+�7M��F8�?�s��!��t��9�Ty|��X4��"��n���X���VUl�r����R��4~5Ԅ�s�j��m���m��B�W�zK�ҝz����R	������
O�Tm �?|NT������9�&k̲G`�='��oqc�X�=�U�yh,4�+	uP%	U0���˝�Yh0��A �\����q�j�>ue��^E]�C�Hr���ͷ%���5Wl�6���u`#�H�A���>R�&�����¹Q�� o!}���S6�G�jN��vD��`���l�!��6�w\���1�����f�DHby"�c��mf(lҹ����aN�!9m��>�Qޭ��䘪��<T���q��@����h�SL3,�ǡ�]��\r�*r>4�a���aH�g�y�Lz*�Ȥ���E �RUUc8Zw����D���i��F��󙒤��)�N���ʆ�~Л;{�dB�*R�	��(��W�2dz�Ƌ�
"�0�t�}q�L�lM^��4}�����p1�./�x���?��n}��>�Y����xR�J��ޞ;�̀JΙgi�
L	$F�mܽ,��y� gj6���G=/��E"��M�%�˅���{��Y��X���-�s�C��?Wb��U������%"qe�x�@��1JvPCI/t�ǭ�uI@��RS�m�1֗�~W�(�ݗ-˟���e?�cwұ��Xd�ä�(��1T����$l	_-G�W�\����Ro�2�����0C�Կ����� e;t�:|$g��A��f�+E�c��Bao4��yae4�&t��<iW������!��?ѭ�jqK��%�3�p�O;�9���������R���q��Χ�5Ug�
{S�!�y�N��(��5��M���dm��D�@uUv���S2u��t�^��1ڲb�t2*��ҁ���.�#�W������e䛍�d�֭�x�6�腡�$ JdD�y5x_:P��A�Ɇʌ�?p����$�`�o|PC�#�5K֫�R�.YoS~�GKq��ʲ��S��dbE�l+^���;Ӌ]���6�6�hW�KiIĆ�SI�0¸
X�7�~���M������<�vu�:��A���T	������K�i�aieT(!��K����<��?VI<�O��G.�/�j�-Kl����E�k������:]XV2P����z]^�����Q����s~U^j�(�٣G>��X��f)imK�ǥ8�([(� �s�oؽ�<���/�n4�ώ+���
ɏ%fn����!},b^=�@0ү�����t�*%��[����XzƜ\i=;�[\R�.c�0�!hQ,c��2�M��n�AByT}�j�0<`��#�<� !�������Y�V豊B�!�4��*w��/QJQ�{�I�̜�?�'��� G2���y��Jʓ�ݲn*��#��U�s���hY�j��'����4�=�`�P��! �v(*!�]��}vR�y
�H���͖��gq�b�!�-���������3/�������B�h.T������~�'�T�"*�!���%-���=�V���!Ԓ*��=��@���C_^���7$�[z�F�B팂M/�V���W>�F��Os�1R�?�Y�{�-,��l�*a	g�L7~�:6�7���@�*�E'Hs�I������&���T����1�F��&	~=���5Jor�rV�����B���uʆ��X6��+����֐fM��Mm����{��t�=04w��i���T Xr�ZD�I��ͥ��=W*\���!�C��l�4�*)u�	�,3����.�����1���:A�Cۢ/'F��;(�E=�9OHX���$��F���F�v�|�P�����:�12=���4aj�$�_y��'Idַ5[$����[*�j��?��>U��uB諔��4C/��Xd53������R�v��p������W�&�]Ե�E�x�����{:	@�=�|)�0�֞���B�˳�׹��#��Z`1�7B7��K���
EGv�@3fx X���Z+N��μv1.|m���G[�!������A%���F:�/� Ȁ�HBʇn$ߥ>�H[lz��X+5�(#�_�fG��R��PN1M�"]
K�IH����o��������P7QuބlB
�p���t�fZ,%��3D'2�Գ�pȈ;�V;K�ዺ.�AQ+2Z�v��k^4�
��� � E�k
���o�]�@�l��n"�2u㥅'�:��ܻ��z��ͨd�F�h/:OwRb"Z���tdwr�6[U����l�H�zy� 
��ӶF��0�, ��Z�#�<dZn�>��j�T%IS>�����{$�P��vٔu'�|�c�/�$���%�fU����R8���pp[|�Ub�\��0��	�^�Q����t$N��1`�o����=��p� ���
��e�