��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_�}ܛ��.��i�F~�~{�J��C�a��K-?�<�>y���yewY�&�_��wr��� jK���w��C�Hxj� ۞�
P�D
��6⼞-E!F8��ؤ�Ct"�<&���J7I��5�@�����-<Ȱ�c#�T�j���Q��X�,.��;3K�_��Mq��.>�V?��Lp-ܘ�jN *�f��7�4>�"� �^��w�i�yG&����a��4���RX	l1䨿;�*޷�}��Ն����.*��`+5�a�u��4j$�[�#vk�~y 7�s�]>�'���>GY��l�]Ry��W^��Ze������� -����={�&`_Ǳ�l���HIS�1�[���u�`�gN���ؔEr��"nU�>E�X�U�4�/��'DeqvMIej�&��;x�$3AJT�y��f,�+�$� �C�c]�Rqpg���O%��0�g[�yÔ�ȱ��D�)�&o���/́� ���0,l*��U��)��=���Q�-�!E��ԝ�b��
�l��j��gÀ9��g����!efq��;nX?
i$w�8o�(��mӨS�U@�7��{�4	�����Z�_X�^S)�u1���(o�v�i��vH�j�7�q�6�<˜\�C��ǂ�x졙�ɶP?�� �r�.���dXFw�� �l�h4������AH�j-�G�kNé�!V<��h{�x�VD�Deak�kyT��_l�啟�Ǌ��N��Wk0�*��}TS����Ҟ��Ӥ ��>Q�tGQt�D�:�T�i;��,YU�/�p���5w
���}�8[��$��Xq�`�s.2����� �Ȕ���&�o�.��3
Q��?s�w��C�"���)�t�!�,�y�`�#_�`)��^�:|�Q  ����M��� �g�u2���[D?��e��8�Ȓ\̚�E����Ͷ�z�[0}��4{��9m�D�-FI�Yk�H�h�2��S�d�;����
X�	!��gʳ����A�[�:�eg���1}6vk�>�v�7��;��p�B�č���f�sC��z�x��$۞v�gA����׋�B͹���Qcm��l��IηAUa&�ЏaF3�N�$ ���̂���3�"�pF���_�]_ī�B8�w�-S�?݀��/ �[�j��T��}��<���Մ�f"��XS8n��oj;���d���<��- k곋wszoe�GV�d�֊����js��DX]`�)Y_�hyd��%� &_�� �
�|F��}��GA�7vwf�g�ֲ���<w�@�R. .$ޒM�e��~Ĺ8� b��I�v	v�+?��0~��)�)%����I���xпJ��QlG;6���qŃn�{�J{�֤��u�:v���D�HV�U�/;�̌����(�*��C�q�t>�,/wО���:eR:�B��6*P�������_uq�		mDz��ei[qŀ/sԵ�@r�x�E�x=����#D���Q
�������‮L��I~�BVv��睐��1��(��2��B`*�Y,�I,-��%^Q����Ŋ2�hB�,��o�+��>.�_�
EO ش�V1���|�ؐɜ�{�er4����`CA�i��ØG��X9������+Br��7V��� x�)JVs[��l����BS4����z��uIW�Ժ٣�WO�u�3P��ɒ{�W��
4�;�lΣ�SZ.l���M �j��s<T܊�t��W�Ǭ�~4�ܯ`�����N��%���zYB�7>�w�g@k`&W���ި.<Z�ۂp�^	*o���9i�d7�X�25UE�~'Nj>�3��@��_�zݣ��z�β�<|P����?�bBsF��d �d�g˞HZ�A�����C�t���e鋍?�c�9��gH0��)**���xF������ȫŧ8{���A\��s7�}�r�4N饴\Ёrǐy~���{�,�g�٬i�a�T�r���qI��~��>Ib^����Gؐ���nO};��[|�dC|	���Q��Ph��@h6�S���$-�/C��Ѹ�����Сá���M!F��H~�����{o^��}z����[�6Evu�4A+��c�D��CH�.����b���!�<�؄�(V>qA��L*��Bg���"7O ނ�e��shO�����b���G�M�Q~ٵ���w�i����1r�1wc�������\���O�~�p��>�%Id�Z>��&�~g�R|���N��3sC���P��՜DDD$Ng���C���C��7M�v��'~�X�{��TlFf��w���BI]�S��q�ƬC,���Ti�TBT0$�ۆ���e��ʽ���s>I����E��Ѫ���/$�Pk��ޓ)Y3���gX/�s����dF�._� ���������R��޵GϺ�[����z%���ݼ�(���9zN���,6^sq�6h�x��0��8t)p[��0��O�7?s�HR^�-}LC_��F=�m���Cr�/��<���%���]F$�=ƞl�M4�Ρ�b����8,j�Y�;C>��DČ� x��o��"=�Q���`B���T]��eÔ�����R��H͠]��3�9Bī�감����������s?�	�������m�x`/RM�AR��o�ch�J�bk����C�����CJ	x&�F��NVT_�Y���6��;j\B��`[���g<��,$W������C�|�q=���갍�s�qc#T��9���e ǯ�Иr%�<�Rڡ������-�!��r���H\+�M�[*��g� �����Cv���G�ƅ��N�R���K���}'X1�� ̺HvV�kfn|�C�dK/�#��_��]9�K���Z��| �{�_D.x�܉�֖�ԭ慔l�$T�6�N�VS�ﻫN&��*��ʻ�P��`��o�㭷�Ց�Ę�"cz	Ժ`f��j/���߄�u�XN���.�����{!5H�bʍ�;���d���9�e�ȟ�R}%�Ը�+xh�^��f4w	�}qg徢�\ӯ��=�Oz�=�HXP�*ᴝ�Q��zS)��A�*�#��`ǻ+����k�s�  �hi3M�̂�hӐ\m�����o�?��J]�{AÐsh�r�-~8�3vB��]T�����8�#Y:B�p#�Oq�X�h�;�7b�H'Fl4��+���q�]����x���������J B�xC`��L�+d��� {]]�D����Lμ��F��Y>��
��7i�"ߏD��)�]nI����`�VE��J]���Wo?���2��k
�ME����~KoNëS:��d)�BN\G�u��g��b�m�� �	~����G�N�,v&O�*��L�0���+]��t���)��!��5�W�C}HH�-�&^�v�u�eE!�껁��M#�;_!����^�Ib����V���O�=q�`�-@*r{R�u�k�O��3RR셇J���l��OoD52�В�'��YĶ0F�.6�^u�����s�}<[M�?g�ڝ�U]�R�Z"�E����vx���f�C\��]R�d8Y/E�f��J�n�e�B�������:��zn� ��q�^w�ʏ�S���gj,������]�"v.}|L:F���e� x��j�7�sʵ��#���]��&�Y��Ϸ�h�M�p�����i�65�i@DJ\���򹅯��_.9� ��̻�B�j�;�n�%r�KpH�\��f���\񊋰÷	IJz��]��qy~Ķ�!�	���+{�����b���m�5�)W��⎴R�x�j:1�D��N����ı¿%	<��@Y"�ހh���؄ծ�DFq̀�W�M'7�q�W��x��I&����Ɂ�MqA��챁R���Åܒ�U!=D�Ǝ�P�ZQ�ݴ�4�;�?���؃Ն�%�hWq��`�g�����q�����n^k��D�o�		�|�k�:� B�!3�+���U�IHH��!�5���K��jXPB	�/���������ߞvV�0���ڽ�l�8Pv�_�X�N�>[�X
��$�%��n�q� �?E�Ѕ��&�08�1|�QZէp���O}�A���v^�t@4�2��	��D����*��/�h�C�����.�P��R��B�6
Q�D�_�jޙ(��?Fv�{��h�2��#�?3(���	 ^��S�UAU1r���ZM��3�80LG��j��m�.�K��|WN�ެ��F���$�]�[�е�#Dg��oM=G�D��c
�M�Y��6�AXz��l�/s7>P���6�ٻ|45e��:b�p%/��pjT;���V��+��i�����5)]B0�Y�?�6p���E�adf���R���HuT��Ν:_s�GD�J����6�b9y\�X-$Ί]Ɍ"����.
��*t��Y�)rTKD��M���B��}l�Uh� K��=��V��
V��&��ް%���X*��Z)���R���PtP��3�?&�
��_��X2J�Ơ�o�+�q�,7r�cU���zع�V�O��d%��p���j�4�9�ӷ&㏚����YAf�ǻ���	�b�|Qh�]�.�S��8`y[֙�/��I����2$�>�B^�j�ć^�Qt�����sm�i�V��1�yh0L�0@K"��j�o/��b�?�rP���3C��b��4e>?u�"�<n5 []'!(= @�Q�H�X�T��XE�ݻ�rj˸N^k!�;�����w^���m9�?�m��棝�Qv� t(�^�a��=�"A,��fMH�'v#���U�j#"�m���W��%����K+Z�}�	j
�����&c;��fj��*��_#�ŞE�@��˴k��_6�@�^)�߫I����V�� ��;麗.�?�0�8K\�8��fc���(7DNn�XZ.̩*�|�Z�.+�k��ą�Oc��)���m���@L��Eam�A�ts�s��.S���[�[��&3���͞&j��=+��R6���� ͹�4فT;���j�����=r�塚ds�j�ݙ°���$m�]�~rb���]����<Y���/���.Z���۰�}�=f�0+m����q�/P^�7�� u��(�/>�rX���O�ͤѭ���5j�hb,i��sb�� ���=Mj:q���I�D�_K*T�6hd�' 2���^W���S��T�bK�s,��f�@Y��G��{�Ͷ���%)U!���M��+�p�YB�u�oM��;��l?3���@��5��hƀ�(ϝ̋��Z%�����;��Y@q}iUP�;����ߍ8d�J���=�Hfxu�S{k��ά!���,�k�*ۊ�|�1��/(J�"�� ��l|Kb�_���}?O!E�zx���4H\1Zƌr0x4A�--�7f|֯󽩞�,`��W����7�XK!�ӛ����F5�;���V5`'��ƚl��!���bQ��X�]���^	�v~�X����w<��h��ڼT$���~��s�h
���[Fs7A�xh.�F��C�w��p6AeD��3�/��ݎ"?s9ՌI<E����@���0t<���gd��IY,S��K�	���r.�����5yxq^"�0ǚ�:bXb%�>�Fh�x�/��<��uf�<���Q�u��+��c���E��j+~a�GO����;
"܇�����1�º��3@C�
,�h����ql�<*}vh������b9b��2�|���/�p̥���rޖ:[���Q2x(P5=�q��K��a��Ȉ��̓B�y����_��CsӁZ�!�;�|���$nQ@��O���,!��%+����d�U�"'���@M������}��7�M;��U.g2�;�y^7�Q������3�ޯ�㪈�����B�|ü��g,��$�Y"������X�F۪�	�{���c4����2(6�/���������C��7��O�YA�j��Is�Da����qr����زF��0�<|�����.&�ܩ�l���Y�bχ����\�\��ڍ�����_Xԑʖ#�ݟ����A��g�{�3��r�F������vj��#��\���7O��F�a���zܧg�K�H���<rLj���ۙ�E������_w.�`�@��?]gS
�1��Y*�SőNU<b���`�CK��ny��c�o���}���#ǝ��Aw�X�#oS�AsUԇh1�ٿ -�*�=�4y�u�\�^s��TT�m|w]�aj��QIn��<�e��K!�\�<gc�N�p=����pl���D�c
E�_���禓�#��������|G0vF�l�c q�	�7�1cfO*��۽z�I%�.��T�~5	Ў�/�JFuK��z�����c�ryu��`m�nUo��ˋئ@F8�W��zQ�&��6�����af�^2�ƀ�d�lx����/(U"JA�;�nQ�H��͞/�[tTyt�&�Cx���o��庱Ռ��h�l���}�����fo�Ao�<�`T�����o�2��$�7�p�W+ A�J@W�?Q�b����m���֣Z�����t_f�0c���w�A�R���{��\�HH�UH�%gh�/*O�M&(���r�2`��3*��dڋ���9�R�39|�{W�t]Sl�\{I;M���j�so7���4˾�h�
�./Sj)[I���U!țд�-���k��4,=�|�b�����
��Dhd�������p(�&b�����LQ�.ɴr3;��G�1�fO�@�K���2[9,�%���������ȮT����}�����ꓛ)]������ڛ;��zY�F� 4e
"]�6 ���\��CW�yy�e��OM��&
�@Ǻ� ���ǻp�|��̲	����
��喂п����W��a�b�!�'?��VE��Zw��}��)b�i�0�v8�<K�y��@�Bܬi���n|mڿ1!����$��f�B'��8¡���|��+ n|+�����3�V'���OSY������P��Ŏ��t��L������!��au�)�(��Ө� 9�>�G�1�Ѿ��E�9�ӲH�;�fu���ˮ)�m ���w���[��g��Bf���8��ҡ4;R���^'�8��A�(u"�����
?$�V�[��+�Y�rtc�d��&��>�a�JK#�\����W�����lى�&��0$��X��EI�S
��C�'���P�7|�F=g>�I��Bs�z"�TRA�sW����9Y��а���F���Z�,��\�����c.q�h�Ԧ��Z�w��4���aR�R����b�L~�1�7�B.�:1l�˴��[y���5w��2̌wʬ�*�}�`3}0��G95���p	<_n;�ƕ�H0��$�����x02�3ݯ�����^_̻��H���PE���oV�A|==�P�<��;���r�Ӛ�����a^��B���mF��E���j?�.!��T2���vVv�i�5��B}]���H�xy��hհ�߼�o�J��i�`�Q��}��g]�}`��,��y����(�17	M�����aȝX�X�$�l�����g<v#�hN'F_�+�sK�e3�΋O���D="�c��Vŏ�r q�Å�bP��pvp�d�Ҳ�I�c'�Ǚ��c�q�a�*`�Z�@�-�t�:��"�+V`�/il@�ʙq���8�7,���@��ώ5����踧C3z �|��n�h�|����=j^��C�J�U�
�r�Ż�
���x�E*���O�z���DO>�K�hO�'�~�ջtʊ��\l����â��Ҍz��
[�8��k�J�e<]��hB��3]�8PZ�쀥��t���Za=X�7���I����{x^�P��T��C�EY��,��"b�i�B�֛f�
�, @���M �B��u�
}������5o��T�a��_˲�34ʹ�8J���wǳ7���)�Ye">N"��|lmos�q�CU�Odl��x��yc�� �����J��Y��(�{T���1�����a�ֈ\&��FuRL}�|�wѢ���Am�����lf�X�	0Y���oD�(Gi�����hXK)(�K.Z���	��{ ��~>ߖX��k��H���D�\5�Hzmi�&�'���fs�I���[���l��w�s��m� �~ע5��vu�!�Z
Ga���^m�鐎���ߞ
�WM3�M�.µ /^������i��/�ߑ��vK��Ud��$�}��P�ܚ��~[�S ��K��A�1�o�;�I	�չa��]K-A&�`�+�?�x�8�,�Z'�F+�LD�E��z};�шT�g����#0�Ж�t,�T&��X�FK���AG���j�����%{mk�x�u�*��{>�L%AQ���v�zԘ�>0._�a,�̪pp}�<'��H�1�jA2��
��+=_&���)g�))6�.���G��5���4�`:<��:�M�O�>��G�V�=��"�MF`���� X���	�sN)b%�qU!�e͇\:��f�$�n� ��k�*\q�恼1���]�D���&o@Ϡ%b+9F��a�I�	�W�T^O{'�0
U��ϩ ��|x�{��ڼ�{Պ�W*�þ�k��	��d��!Ҧ{�@t�n2)��΢��;�+�S��#Jy��a��{�����[1�q1��3oqvRac����+�X8�5 �_ƒ`�J]fj���%I!�1A�s˺�1�l{��x�e�<�e\��N��Z��,��S�K�.L>�Cp�3]�x!�7ħ>&k�N�
����x���֏���5���8\�O֭dY�u�e!�/�V&���4���F�d׺�����2Gz�g���F��9�o����3��[hZ]B@�.��NSs��w�u���%M�	Y6����V�)9�Il�*��q�R{˿j����~�� xixJ�Y@�O�&$��6,�VW�̰\���W��2a��mꚁ�����������LĮYy^<�n��^݇=尪I��BlW�v~_Ns����?��K�*P�WT�p����� ʏ�-�X�">́|a!>\��	�CNjR��ځS�����7̚[ɸ��ѿ�T�6�|����-�B���ȴ��piT�:փ��A
��
��o���R���v�����ފ�ԾCտ��h���������ȷ|�f�/�EP�+�QA�(p���-�qd0Oq ���D�1���^mT�d?a:\ٜ�Ε_�M�t�!�o���S�e@��pH�������������cw�˗�h>�Z���������N����
8!��yRƌ���^!2�~���8l����B�B'��Z��";���!�?�?�`��0��b#���vRg��kM���%�2WX�1��:aF%�t�� _VQaU|@�U��A��(& �
a̘�խd�s�Z�>��-tQ�kB�$����gExx��E�(!�'Q��H�����A(���]n�)�EŁ�&4�ha���^Fm�>�]�%��]��B5IBb*��1�&��Ԝ\�po.�a�J!6�}�gBl�K ��D��90IJ�:5�E}�\6��1���� vڐv$/ׂw-�ο�E_>�g� ���.E�{>Oj'�	��D��j���s���"�F����_)�O���m����Sb�2�Н�eUq[�D�!*P�L��D�|�m���CS�*��+�����c΃T�XU���3�Y�Ѩ8�V�%(~��&]e׷�*�IVgiyY��\�����M���O��y)���o��?�x���z�G�S��;J������EJF���A!E����}+3S�@��k:�	r�9��2�����z��KXS){�'�i��J�P)N����ԹǠ^ʮ�V����y�˗��hY���x��Hd;/u�����L]��%A���l�ݿW�I$t^�3�a��$�&?뀕$�m�@�L���%�{y���K�þr��Џ���9'd����}@�㾳���V �	�{J�C����b���K�5���L���掙]A]8�#]�]�6K]Є �ŇR�X�/�?at
���"�s���hʑ	���(�|�ר㛕A��}S��JV7O�jŰ{��W<=k=��h|�0��"IK�ΕC�23�����\£ݤt[��a7�O!<] �t�{؊�7��"U�8�.�5��<���VW/������S�1�L���G����Q�*a9��O�Ǖ����`��V;��/���X�m(�>!��phl�:}��c��۝����p��\�.��B"	3�h(�M�I0��;��b1Cy4����;���V!1jCq��At�9yf�Ơ�%ؾ��'�0aD�R$���`{,V�����%����ֈ8�R_얁�����j�v�)^�%�(3�Ӧ�����3�-���,����T�8� $>R���G�5<�?
�e����f��=��ܳD��xXh�Y��z����?�U"��I��w��3?X��P�S	�1�AW��Q3V��Y�O
�,�Tw��޹R�C�@8.��х�6��]�(���<�+�r���vǭVD��\Wwq{�ϰ���R�@�H�n搜�-.�Y�^X'٪b4�>�m�s8�����'�A?e��WgW�¢U��˻�[?E���.��(�;���((I1��~,��w8 q�fR0�v
��a�8�EД�}���[�d��V6��C�[h<ҥ��x�vt�_Ш�+�k?�Ŝ2�tyV��>_���lx�%t?	'�>z+��&/��*������s[���W%���6�l<%9Ȇ97袧�VQ�}yJ����~ ACf�ӇvB���wYWKP')H���q��ڮ7�(�.�x��=L����2L)�O���;�.��;��Y��`���EyIP����#��� 
���]1��SRZ���`��h��)(��
YZ��e@���c�ajo�ڱ���
���]�~J����Zvp;M��?w�0�@�b�V���nh��k���0�q���q��/��*)1
���F7�/��":�D �۟���B���,6v��R������w��X��ʖ�V��	��-�F+MCV
��X��O��\a�%'y�����s�����pW��Mfgk'j���;�"]4ٲ��	��bds�?�A�/�Ę�݌�߬���l�P��z�A��(J%�fѡ��?/��B�|A��8�9oF�6���8o����d��L,�r� �Q�j֠Jt��B�̷���-���f!�B�P�ӗ�9
'G!��$3��C� ê�WkN�:fչ�p�[(�Qn�^H�>ˮI̳ʆ���F	#n���ؘ���=��fM@E��;����K=�f�+��ҠK<�|xI��4[�N���%u�!c�̰уą��V��4M�Q��������S*?��W�j-h�e�o>�_T��I:��Т�=q3�Ȗf��{���2���)�Ȭ+���JxK���up���������l-��cF�������8a���q23*&�ԣT�y��pd�@�iqπީ[�ҤG`dR9�Y�8�^`G&Z����jY�Ӯ/U"������H^���r�����&C����x���#���l�ՠ/�v�'.=�yR��Klb�wb�T�բl/+�¶e� ����v 1��w���%�k����/Y�R��%�a�eP�;�cB6_D�?O��oB|��|8�0����K��r)�!�����]Ԓ{ =����[`�F�� �Ơj�L���|&%���;5��3M7`�8�u����g��^:���%A�h�7q�'��|	�i)x�^i�Ttc��0��Zjc��P`�����~C��=B���,��ڨ�b�8����W��((����n�
��4ܵ%dV��w$C��s�����1o{sJZ6���ɖ����r���e��Lb>�����Ẑ�g�W��!���t��Q�|s�Z�3��r�G� �@O�L��P��5M[�\�E�hP�cP0lwsJQO "��E�*	�e��m:_����xH�v��r�_�j ����|�����]�"�Lp����{�˦x�[Ԅ�ߗЦ��o�")��~��$�
ҭ�;�jrNg��2�kD	��bq���#냪x�� ���K��[Wo��L��X}��W����l�y0=��xx��두#X��dC�H�bk�Kȱ<B)ԥ�E�0�m�Jp�6��C�z-�Y�qn�˫E���<�%��7�Cz����҇��1S�L���#�^a'�.�g���K�9��Epz:���?���Wb��(n,K��.)��TFIn`��@+x�/=H�6�m�*����.[qЃ�о�ʊ�$���y��>��Ӻ��L�q�ю<���F!���$�(Z�Dar�����ڐ�>�9�(\�A�T���Rx?�='b��~ȷGk���_7�[�|����0�&��렾:��;<��Kj��Z�T�0��n"��:-ݪ����S�2� �&��2��ս���θ�d!��mh����8��O���˚���y�{���B���b�s7��ȟo'�����a�J�L���E�	4k�x������ʑ��z��r(F:����֦pȫa4wb\w$�=S�7yͬ�f ��������_��:�H���C��M=i,%a�IX�+1�ዲ&��.i��S��P8d��f�1�+�T��'eH�mOƚ��jI�'��ܖ�]�\T�ME������uF���DtY�l�㿀TiVN�.	|4qǉ0�bC���y
��77���+�������߃�S��ؔ�s^�C Q�8 M�����QtD��L=#��X!�#.:Ԃ��x˵p �8,kDYI�m"��)�:��D:����5$ ��2s��5��ij����0����=��k*7��D�d����U˨�cD��s�Mо�4i��M�� �5��?��~�P(�L�JG��q����.� WW�J FS4G���֌���S��x�~d�7"6�g�ʓ79�i�r�>EhbՆ��@g�����JP϶$k��o�E����/�`k����o��!��/�&����bij�-o�q1�>�Sg�b���+�GL��)�Vg���nҞz�Ȫ����B�6�ht��O8I�v��B�DC����7����#�R�젛T&�"W��0�8��������^V��gD�6��˿���P_m�>��0=�c�q���_��'������ۍ8{�X��oS�o ���L��T�נ9��)�iS�y���e�r��+�x�C���-��>�V�Dw�j�O%*�i⌄�T������o�U�[���"���]�f��rm�4���y��W-Z[%��Nf�~u��L������g:�05C��2X��Rd|�N0�Pc���8$�Bj���@��V�ڸ���P[���7<0d��FFݫ�h�r���$���"`IK����d��ǯ��mc	 ��S:I�x�+��'���lj�f>�1�� y���䟱�5�\�#o/��zq��ʂ͗�D��^S<S������{�p��p��h��{��c�|�ݿ��*���PI�E���j�j��0Lϫ��ݖ�i�X����8܉o1�e[TQ��B���B����k={��`�̜�V����Li��#�o`7����-�c�-��f�B�V �&�S}��$�ݷ��QS�&܆���ߝNhV���;5{x�օ	.�5�n�m#^�}Q�C�/�j�����;��C�F��{�[|��_]�P�Veh��1
W�����W\���+,8�Nt�w-S�N����w�0Y������p1����\� =��BM�n�-<EI̯R����`t�&y/])�2�՘L�T�hrs�d����15���۞�:�[��Q�pn�\�?��[�g�1��Q�$��Ѡd���Z5}\�mr��F�h�4�y�O%�9)�� �֙`t���K\��XtX�oe�(t⷟�a�S��7��{���ޕ%��@ʆ�A�~�U�,d+~T���?k����琭e[L�@>?~��>+g;���{F7]��e�e�@x�9�������\I�Գ���SV��i ��G(�EO��"�=s�di��?]!�~��xl˕zoy�y{��a���7㢓�|������mO�kX�$
|��s)Rr{�gz����_�F�Qc��)fwM�P�!��@c�jbH�ìd1�1�����}e��I����;�h���3��z-��2�
����Y�Z�~ !Hn�~%#MRnl������O8�G�uOW"k��-M��XCE��ѼVj��y���yح/~�0��o��v=i��NJ���&7�v!͞|~C�2��QF1�M+)�R
��[lau�l����xO�)�F�����\X���x��.�����b�[؟�jߘ��&����ϊ"����T�}��Ql"y�����Ƃal}���1�c3g{��r]ҜL)�ʜ��Y<c�Z�V�}���t��]0���a�{���)�)[I�H�E���Μ&��r��]��3Z��Kt��V�V#¥8����i,.i�8A�"��=���s�@Y�oe�2�M����VUY!|�_[v$R�'s�����6���ve�2��>$.�����(��#>������1*����ջ5 F��Ȳ�@�Nw�]�̙|M�B��ӑ�pB=�V�Q��+�i����`�_v}�]�~V�n�¼��Ԡ�0� ��G�l��cI{[�!���#����3��)�cU��)mG���2m������葐��7�P^��cf~�TZ	_�uؐ~x�$��%"�[5�vimbQO4.2S���YR�
�'(������o����2��"�N�kw���Uh0;c�]�[�Z�����dv���;6�.�lE�yP(W{B>������׃�^��ǭs��y�(��U0�ЃMjn��N����`�1�X|_�]ܭk��K��S��_(ݦ�Bp�>��H+����%���Ҹ:����Y��{n���F:ri����n��y-��;)9��X�����:��B��`6P��������M��$~����x�3�4�I��3��tZ��"w׶3��Q��5�y[_��w&J��h\.hJK�D��ĕ���gI7�B�،�� ��
��Lŀ1��UW4�������Y��m�M�̻ípv��2
U<�~���JY�p�q e}cW58@}��4m�DM[C>�Q>�/����9���o�.ۼ'��]��f�x���͜Pp���(m��H�����T/�92�ɚ7������#Ǉ#�2N�uڋ+�r��p�a�n�3 ��ܘD���p�	�� ��C�6S;�%�r�X�v��V��B�~Wܴ� n��DH���e)1��/�&�)xy�*.�������oW6�4x��(��
�(ؼ^����U�c�!�i=�{�����4���].�Y=�Lۘf��wJ�5�(���	�C`rm��Dd�e�=�>�L�m	͗�)S�����pȖ�^3J �g �F�7Va�����ȧf�Ad�2�=Jz���qϵ5�η�`(��X�S#�^��jӳ��,B5��v�4�-��QJk�y���������
^���`V�����x�Ap�V���n48s���]6���x�6�W1��!�i��E��V<� U�Z8d�1��<��K�J�I�m�"�l`\�?�0�q!N�wn �~�̉F�
��K�5��r�L�KV~�n%��"u���[�N�L2�if�������D��պra2���#@�i�J&C������	�䷁�VLs�k!�"�N�r�e�_m���SV@v���*.=օf�>i%N���G�����g���,Š`�Nu�����S=Z}�Q�0nF���$9��w;�m���r�Ct�]ѺY=G�=	���$�`�G���J����X+�}u��҃T��t���Z�Mbm�qE�0z{sw|�9>��8�Ex�J���������-PP���<�G���hk��y}|t4��+W+�rCҚ �9Q����U^+��枿�c���ۡX�}���\�!��C���i!J@AJ���b�kDv��x**0|�]3�~bP�8�!�]�b���1��Kȩn��qM���=�uC��#�>�Rsm�x!�v�`�i�b�`�?�龃�����c��#v|�F��Z���7Rx�3u�6]��/�"S5�ׂ�\ϑ���Vc�J�eF����c�Qc~ ��k/�����rTk�m% �`ܜ��*C@�U@�w4����xk^�Q�`�����IO{��^�< �@\fsU}n��Q��7_��+c�M��t*E���Iq��� )Q~:\N�D-H/ak�]��urL���3;��;CA�κ��vH��=/����DSJ�'���^�b<�%��L��/�nnl����8U���,T�������9�m�P�<x�Q�#��*�𚌶'�7��[p��_IH��	��ܢb"�����)_��f���]0Z�ҍ�m�j�X�����Z�����g��h��tM	����a��|
j�z�d�Oo�R��I�ܧ��P_\�kw��I��FD�e���̸꣊.Y`��tk_���3��++��$�\48j�!E�S�u(g�h.n�l��n-�_~�u�>T�/�;�X�d6���-bsO��$M=�f\QB㌠R��i�e�C��uG_۫T8Ԫ#�\��>?��Zt���S�˴-|$����:�U�࡟ OMK�v��
�h0֝���:m�B�x�=:��ܠG$F�:�� ��gyb  �k�чY@1�{-�9>xt_���\��Aa+�d	:RX����u�Ҫ�yi���I�̝�˜?Oi����vde���nd�7�&�v��2Y�Rk�'�r#M k��gB7���{�?���MXB�.�]��yGÔ�{������T��Hzp�=j:t��#;�I{�v�^]M��;��1���--2��vw��?vؑ���+p�AR��Q)VuXk%�f�2��3nƑ�Cn�����U־A�v>�x�M�M��Q�;�|�V�ev���Yb���ǀ�6=���Ky1���kR�j�<�*�v�)��G�`���n�7f�A�s={��h��쓼e�ٟ��u�?�Ę�W���)u�֟����p%ٖ��do1�M�������R\�A�:���r���x�]��خ�#.ٲnOɵ19�v/��, �:7b��i�������C���8�3MpXZ�S�!����1�#'����Q���s]fQg%�~ͷ�L*������%��Vŭ7��cT'l�B0���b�~<��14�X��� �MfM���S�)B��n,�(�u��1���M�j��/�w�Ԏ�]j��l��?��d�x�#���NY-{aN̻�tNέ/<l�CFAy_���)��v��y��J����V|��1!�%m�K�JF�)�X/�n<�Ơ
�#$�IJ���X�mb�`'n�P�y�koK٨0�"I��$�'+���T�y=��H>2}�<�foC�V�;}}ْ� ���,�jR�w�-��/�VΑ\����[��wA� #�;����K�<z$j�x,��t��pY�]�_�h�G^�H�lP����f5�sv�����u/Ϻ`�geR�%R���p�QgB��v���w5��R���΃���j��������}o5��ϳ*w(����-v�Nj�?�{l�� ��[�9n�TO��� (����������-��+���AI�+>��?��B�/Ի�ϘI~�4c$�{b����V����}�04��T�\�u�����=�<A	e����_���TG��-�
Fh��DeY�����j�I1T'u� �^�A�Sse'�K{}�~��}�r-2�GZ��,��)b!��_�3�]WM.q���#�Q��xE�	]f�����9�WkK�Q�i��E�->@��PF.1��n`�у@̼�T�=�a�U �s�M枵D�e}��D,}��8���}&�E0ߔy^#{u���ځU���o�9���B���ގ-���Ks��7k8�b�����&����K�5@cCapKo�
{�`Xaܝ�[��`Dث'�Rj�hII"��&���c(K�ǃJ_sE�1��O��}OH��B���X����͐T�rA���:A����~uާ`��- gj*x�Wn،Ĺ�)�>�~fE;"�*�o��Zx	y�j�v���y�
�19��K��;�%X��0�{���u��'"��J�G����U���v��V�g$�h��~l.a�:�F�ε���M@�8�@������Ӽ:)�?�L�C�#�)SK=�'n��'b�_����}{޹�W5�2c�GR *����v~W���[߱�i�^�\[K�
��!�)��R�Ѹ?�i)@����ag~�X�H�}_=�d�Ha6�7�Q�s��3�&�C��� ���0O(�*�t�����'s`h=Zӕ��-�l�F�����4S��2�3 ]!An5��n����uX���A�/�� O��o�g���F�����@��)���dX��1)��H��fܥ5��L���H9�ܕ.]���l#���!�=�-�x#���n�4�����N��o���A�K��:�,���zp�G;_��S� _�+`�B�ĕB�Y [��Z�O���9����blf{���d��؄%�|bӵ�A@MƠf��vj�]R���u��0\�1)��G}�u���L&������ �)������x&�y3P
=�o�z��B!�Yq2�a��_�v�c*w73L:�S�u��3��;G4XS�%����p ����'�v�Y�(��ۍ㽤5��������_�݊�c���O����/�F%:TA����Lr�l|&�p�F���#*�C�>�9�3�����o��<ͥ�l@�� F�1��{Zޅ����=ue�������=$R6�*�WIȟP��E��V��^���`e�l��$L�)�ף"�/��o��P��3�ٔ)���lB���f�Ҷ��r~t���Af�I�ʮ��am�}�����/x���P N�-�m�9�:���.�(��(ߊ��r�?����G�t4�A�����s��md������&����ľR����K�4�Y��.l]X��=��$�]����}]�9����<r��JUHJ�(��0�\��=�Y����r�9Z��T��f h����2	8+��E�8ؔ�Gxd�uS�8�������F�gqԧU�$�u�jXԵ{ 3�um�Zϔ��߶s��e��h������v+�x�Z�|��}׳n曬���
1^V
����|.uZ��{��� k�eN���(ۋiX�"Vu�E%(#���U&o�W=��nUU	�������0���6졪X��I�m�[j������#2O���A �/��)�L=+��؜�~��)kٍN.s�#*	��8?x�,xʖ��"Cٱ���M���=�C�:��h[�/?]����m�[�e��׸�*���B.
��;��w�G��sb�2! �u�w�є�����Y}R�߲�"?K�Մ0��o�:�W�3����\K���X��}����gP����"z"�������L|Xq��"Wk�^�f:��� �[��h�N�m¸�
�6{�c��܃z���
� j�G41K�����Z�l��L�K ������ׁ��,%��h����
f�R% ���+ɾ?��������_q=��/�sv���py�\֨��@L�5Fe�K9^J���,ED�d+��p�R�k�OhO��Z&	�N]�L�|R�N,6&'��h���F���}e	�,�1�P*�Uh��E�ݿ��f������‍t�Y��p���f�X$���.eķ]г��[(ǹ�P�����=j��ݨ�,�����u<���!�Ϭ:ܐOʰU�E7j���lI�X3���ʠ�������Tg$���)���y,���cz*9���a_MdM����%<V2݄�i:uN�q�W�ؐ,?�`�`���\�b���|F�$�V,�Y�Ξ����Ӑ'�:��v�嶠Wizj@�<q;H,��/v�	����y��G�7��2���f�,0�P���k��Qh2�8@�i	%��eL�4` O3
=@�Di���o�,�Y��սi'���_�0�����hR	�5���:|.�iZ�Y��j1�U�$�7���ƾ{l]f��Z�bg~Jcs���
 O�?��L]F���^���[���hi�<DN���i	��W����O�c�WÜ��Z.�OHou�|���;��ǌ�^��SpZŃ����孻X�4B�e�g=���7v��u��tI��?L�P���)�@��b�2�b�ċ�/`n�"�j�T}a+�^c�����N&�]�!��~��a/�m���ü�p�m������(� ����N����l����7<���J�P;l7�Ĭ���"al(�n*��~��~����v/���^�c���$��" ��h����e!T�V ��U��&�qi[��Uto3e�@ǷL��u�3[�P�VtE��6�r��ЃI���̗�rf��� ����o�Iӟ55� �����\fЌ�5m�xe_��E�D�����"SLUi��&������ �>�G(�����-|�<:i�A��Eۏ;h�x���F<������|Ks����<�6?懠�]y����4�f�ޘ���k�h�u��bٱ����vGR��>�ħ�Q�F�)M�]�?S�`�;�P��Ϸ/=�� ���>5&�ߙ��hIN�~T��HA���-3����$�Z2Z��K��u�хi�y$<��]yٗ�n�ӏ;����Ė^}ǒ�B�tN�b�2Y�,�7ã��ꒆ7��^Qz�l�6l�">�F��7�"��ff�"���A�Y�N��[�޲�z�k���୔�K�eU���h^1�-WM|H�zX��ؕ��v��{�0~����:j�f<�+��<�C�r��:@����]]���ڜE���֤ߦ)����&�~�a�Y�A��]�}-�`C��m���I����[4�U�)�YY�]�9�<�K�Y���|:����.0 �p0��Q�P=6�����d�� ���f�??�/h�G�2:w`M�O��mq*랟�r�竲b���ms��\$6��s��8�	���M^���b�|�,J2��ֿy���S�\��Խ�9��F�y���L��4�baO�L;��i͗N�)��pl��בL�*�� �7���R��8�[,�jn�'�N�-p�aⰙ��U`^�֪R":Ǖ3��?�Y4��V��S�8���}��l�,T�����Z��b��?��,jiDME}�&a�U�������X���@ �<�U�5�R<m����gt�4��m�tP�0�@<��f���T����M T6���hڦ��?RիA��hwt��,y�\�t��]��K�Իz�O�
�a��dy�L~2�N�W��f%#�քG���D���|�z��K�� ��/>XFj�k��&�=H��]��Ц�B$:�%�šU���Pw�>���b��.9û�k\vtե�B�= �'r�Q!t�X�o$�zE�U��|o'=��@URJ���e�?$����n 8�}鸉������T�碕�Т3��MV�ƶ[���'$bT|�I��ޗh�*�W���uVM�ґ2b�[K�D�m�O�T�Ⱦ���[9E�*���۝{��������d��Ͽ�P��
c{�U ,���瘻\Ig�>a�~SXz�TO�Y�O�v>�}n����H��4�$�"+me�*9H2lu�)7ţ5D�A�����p�]*"�k��,�H��F(T�:�Lx;PK��-��y�C9ox�2:�L�����T^$X�sAr%;?��c�+N���W�[%�y:滢77�<CM�^�A����q�0!��=�
%+��'�&H�HW+N�D���gY\y�Z5䃡�e��ŬW�o��t!W�͌qF��wB%�^x<�W��_���Q�94-��:2�v،�%�W��Qc��{k�G���J�t���#�����@�cm�[��Y7����	���A~RA�?R�XІ���翿�6�L�5��6L�i�8�ۢ��j��xu*���ĐQ|Ձb�!,�:M�����'#��)مLםiX9�^>�0x.��/G�b{B�~�����z�h� ~�=A�@&�|x8�JC7���1�C�Ma>�?�w�����$�9�̲���,�x7�ȌQ폸���Z 4xMFPr H�<:챨Mlے�;�����wr�4�HSh�`��t������s�/uN´>V/�Usuާ6Q^�����yb�����6�A% G�.ne�u���P^{N�V�V�uȊ��+8a=��b�j{J�������Ӿ�P�&�R�o���?��V�Ѳ�e���vF��=;���C_��M��h?Nv�*L�$x]��R���ecz�r��e%  M��<y
��M�y%�������md�i�Tn�(ms��B�l����r05�.����꿡��˵UF�щ[��>����փ�	�a�2�z*/�e�Hhc���z�I�ܝ&BB�=�񒘛�[,������I�DA�jDHR���I�O	���Ct��\�O�}�T;fJ�{�C��n�}s�`�u�?(�G�=T��������ڕ�{9�f�:����j�{v������}�b`	Y�V�o���˷) �����:��t�K�µ���S`���:L��e�������sE����Um~6��?m�l��Z:����'����vҁ>��%��C��,k��d����-�hu]�+�e=�����;Q|q"(�0j3�$ҿ��~�n��x��W�R�u���&s	��=�B7�_tWD	P�b��'v��W`Zaua�����(��	�b�$�FU�년�)��k�e:� �=��iyod��M"�-�`����l����k�/T�����'n0����v�zI �~���֓��޼s��5�GI[e��G�[Qj�V#�,q����b�] ��z�?��?�J�����<F`Qn{}�!=g���U&��AY	�:���,�|'��i|��X��{0�wd탧�Ɵ�V���՜�V;���.m�DIsr�l��BG�"?���k�Qڮ(	�Ȋ��1ޱ��D=.�~`�vb_�nT6�+=�gub�@}���-B)L��h���Ӄ�=����e�u{�f�S��E��
����(�h��֑�\ =�nu^=��>�v����j]��a�3�/�ݵ��9ƶeop�(a��Fp�f0[<,"��6OЛ_�]�s�wڠ�� 6��B�h����1�Is.��G���e�[q��9�E)̓�����*�c$��J}/vqcL&&O���os��[R�����t��1���(+4� ��ŕUUS��+t0u���DI	ϙ�B�ɀ��2C)��g/.~I��y�;�T���pJ/H*�|C��O���=����E�nIY����!#[��:��T������XH֧̈2�z��߸G���ˢ�5Hܫ����9�5X��m%`���ej~����OL4��jA7�/.�Ni��S��"yE������Udj	'8$w�n�;C�D�-��mQ!�0f���i$q�`��2���p���[Q��g��̋��%��m����E�L�?1kIQ\;��OԽ�q�k��Z��{�*��<�4sc��~�ݾ�x��A�Ӊ~+p�BI�X�!]�+�+��,�����*�����"b{q��}\WL�bP8x�Ad���:�j�h�^��m⹘Ƴ�r+^�Z���!�_��V���`����y��%� U���'0���m��Z����a���Q�\�)��F��=����e�t:�+�-��$X�"����,Dܳ�m	�	���ۤ�V�(�S���CPP�T��ͧ�3#)�D�l�ꛭg	=!��؏nF�ۧ�8��`.9�5<�s}������ިd+ku����nۨE�S���ZG�b?ggb��+�pH����������J�->���Q�����m0�b��K�X_�&	i�5���C���&N_����Gx�f��
���O�0�@{]+�����)������sbX�2.vβK��k��y����9�3ڶ�>zl��5c�&ҙ?$(��[cmza�p���-���8q��T=$�W
��7獄Ji D�W�X�|b
_8#x׸tƱގ�l�FU���)�1t��6�<e:� �������֒���iD.��"8��Iz��5�'�Y��dQ/t�,��:�����r�k��M=YC�i�=��8ɧg��6Ke;��!��z5�>���HsM�R�ϓ���?ˆ��@�l%Rѣ1%�f��Q��9Ц�S����Gr2��C�y7���;�U`�3rо�c6�^ħ}��-��-����M*�d�������8!T΍��n�-q�r��6��0J�#rI��]�^�!�&D�[�4$/�������l���S&B����h)���1���g;���Ȧ �}�/l�����f$8�co���S�F���q��=���C����|��݇L���^�ҳ��\�l?#kI��7�%�d̠tqv���| %�etuU�vf�)؞w&���E�Kp�6�xV�$�i�os��"i�Z'qU�D�e�G�I�Uk�����a�3�=���{�굎�6Z+����԰���ۀ�?�>K�S��S�� L�	���/�/V�)۱
��vu>j�HJ���@]�s�f�T8+�=���[}L	$�� �� ��Jm}�_�����3�,R�dA��/�x���9i��Sb�x��{"�H�eƑ�	/f�M'ٺr ҰL�=��v�����F(2�Z@��b�>��;Ŧ�
̣4)���o�(�Jp1�AXA�dYL�c�0c�O�l0�R6>�*@0n�"^)�#�s��e�c9�znb��<Qx�U�,�lQ�ᆂ� ?3�+y�L�Y\�|.��=�f����1`�$ebh�B�~7A��f�,�u�TL{כ}�z*�R�]����j���z�4����jJ2�;����X��M�F��O���Q����8��XD$��a;��{g͵�c��V�{<|���%G�g�����%�����-)�a&R�m��{����m�X�H�<H/�iR�/�-k-mM�>���P�P8�+�ѳ��
�y}�f��S�|�9�t��Ѽ�֧��t���Sv�P	�J�3���Am�׀��x?"�Q�_i�9��	�Rn0��<��{�mo�<��A�jѬ�sH��Cb�Yb�G����.ڬ���Q��?�璏�\z&g���#���-;�