��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ`T�}�w7�ɴ��劂�;0I�`��=�ùJ��o����grB�K�2�Z�P����ko]bn�E�[�+���d���V^�~
/�t�fdA���	� խ�0~sߦ3)�\��wJ_��1���puMTO�oM�����K��XS4$�
���@����%�%B��f�[���7
��;��~'݃B���L�>h^X���X��F�Q��\��6�n4&+�Ms�^`2��k
fZ��n��V �3�Z:<RNau�l�	�HF"o]���l�����?�Ԑ/d�!e��51/�Ȗo����GoO��^�'����=�l�ls�ޱ�	d8� �s/l�����ZM՞J���H�Y���&$�[Tr�x��S��M���rR��e$�H����)�aVs�+�IՈ�W\@�D�Ȇ韪,�0��F��,Kbo>�}��Aݫ�t��P�Q���c���%$ۏ�(B���>��3�\��P@�IjzA,�oă2t�L��[*'���H�kfo\��A9N���f�%�Fnr�Z����[�JQ�/�<N�@�%M�O�	�?()�$��`{|<�j�j/Z���%[���P�HԼ�u���� vXn6�</&������a��U1iZa��F�V�q��H���d�89#q/��;�Fc����c�(������S��AO��Z �t�d/���&ˋ
ޠ��F_��Obg�Cd[�'O�δ�\S����:�S}�	<Z��#�8*����҇WiG|L,�&?��J/h sq�j s��I�e 60�DOx�M�W�m�ɩ̬�|B�o$nf�i8�r�P�ҥ+?��c�-�̎��0l��ۭ��\C8����8 ^�k��R�$nТT����C۠�?�hۻ��j6i�[P��;4ъ�t�8��� Ys	!���ne0I�֫�p��7�����ZE�v�ƭ��KkB����}@|��\�?��������Yg�� ۇ&-�����,Ą�4�'p��_�4��ji�>gH�����8�/7�N��i���?W�'�)���(�@b��Nd��1�֞J�VH��oⲻ��Ô;�02������:��!�d�]?0�Ip����^�>�!zuw���(�FWG����A�x-S��1�!���>MVs��ˢ6Ք��H� ��צ�� �T,]�Z����+����]��G�ʡ�w��bxe��,�����<R�苀By�����z5B�<DzQ�Pdܲ�>#�h���Vy�T��u/)jN$�����v�ț@�>��7��e�����H�����U�!��ֵ��^u� ���1�v��R�P�*E����V,��V4p��"�k�0��UxG�Hp`�ZcHJY(�i��4u��G���-�&8��J�^�y&6�'���?���7�G���6�f���_�(5��n�	1e�2��q�Î�����,�?Ȥºٍ*g>�'@mA˛0M����w� ff�� ��<n@���Ť�v��6��� hk+��a�s�	J*�0�U����,�"yL��'e�Q�q ��h�������"˰Z�]5O�q�;���l���$�4�}���5M����`U�~�C��r�;��ЀtyOcQ����	B��:|>vڊ�S��;u������!��F��_
�8��w�\6�`�"�Cv��,<<�/�Of02���hђ����(�=y�P��������A��FQ�	�H+{����j,���6X�}�J�5��Bh���G�����T�'����?o��Ԟ�M\�""Ky�؁l_��%�ٰ���&s�,�>�}��Y+a8�]��rC�;!��ոYYB�%�B=�B�L�O8N<�>R�����W�.s�T��@��r���b�a����W���I�%K\r���'9�}+������l�,b��ӹ-��?�c��tB{%��o�vA�aMl�ʽ��jG䷱�0 �~k�R��)�.��X�Ž	S��v��T��/4� t�q���ŧ��L�9R� �3��'a��T7��^��{7+�E M&�<�W̉<,B���p9����sf����9�֩jM8K[F��@�}|瑈���Ypө�'3hL�mR�h\f���I0^�0�m��8Lb甽��(�7k�y�Sg>��w��n-�.��ēU�`髆��]Զ�e�r>������P���$<w.�;�:����ym��z4L��Ȉ!�Ij
��̄��^����u���{��Ϳl����(�0��x�6�����`���
_�ϦYA��ܹn�WW$Z���+�ƪ�<�E�w>�C�T��hI9ޖ�2[�<ry7'5<�x֖��eP���a�����<x���Z6�S@�T8�Am�ѣ��CW�}qja1��Kę���/'��rl�G������*�3Ou �������Q�[lc�����-�0m�ʟ��}R�Ifv�]���x��E�0�%Rĵ;}"Qv�u�f�NH�HV���o�i������SI+���L۪��͸����^)R��j퇈���@�](7�Cyu�񰣇�.zҢQM�hv^e��=���"��	v!�+�F��d�����8������&=���v�̓;]���.p����׷��E���9�0���p�g(s���-��.XI��r`[�Ã?]�Vt0K���v���j��h�kW�?�U�_�P�`q�ix�$�y���JW.�o(x����5���y�����8t �L(A&`�b�Nz��J���2i���jK�hL�j]���j�)6o.Fl�>m�D�L�܂�j���g���^�=O�ֻ&�eǕ�ʾQ"ޛF��2��L��"8��#�c�؝ŝ�Gҽ%^���\����cV������r������2V�ܰWnNY�5PF')͊ ؇~P���3u�u�wsb��]�Qi�Gq����\������j��^V�{���H/r�tƶP��0{|8��.Lu�mr$m.o8�+T�J8�Uɑ��\O�Z�a�LQ:�p,������xR]�Ǒ�0�sY	D�r�'>�a8�}AN���)ǅ諑K<�J"x�"��
�m�J䫓[s�#_k��`�ӫ����3K@�kb�"��Fj�S/kE^�8��6'�"O_��{��EO���%�]k$��	ǈCZ�Zπf��tӰ�T��Dl&�C,P�]�#����.��ަ=g��V��@C)/l=A�<����D��W��:��ѫ���6��E�� �z���q�*�ɯ:����'q�*����H�ӆ�����p��e���ry$ ��&�(l��{q�٫�b�l�,�ù#J��jT���6���R�!�p�p%��6��G����	��"wg�9;�j\��3��P�����،���B.��#��x_J�����o�"�0Qad��� �Gψ�� �'�� :&�qnT4v��bj4'3�K~�7f�����5WG�ؓ*(�f�V�d�H���]Km��	�w����Sf�N�������.�_4����D������b)�{D7]4!_��	c�m{n&;���x�)7-���Ϋ�4�n�0�X6��~d?B�Eɉf{_0���+���mKӰ���o�#�������%��;c]�&BiZgj�F>�_��y">�K�����2C(��,�mǺd�E��ӛ�̫U��o'�s?S�����¤Wj@�m��b��Mc���NU�@����<8�_=0fn����lC�B�-.���K�i������>�ٖ�5�"8O̡��LU
���/s][� (5%��+{d>PK�8>����)�e����J��J(�6/�O�>�E֋���aB�Ғ�ܑ��_��#n=�������[ ~�����6��*���r&�㞿<MU!� .�C�=�����=`�P��P�&�)��3��s����\``�y��"4�.6�E߭��r�]^���r�a��� '�:���;��3���%VGe�4^j���?��������mQlLOB�
�^�������gib,"u%�i�|��G��w�S^�q��5#:�M*�q;�#7 3�b�(�ޟ&*V#d$+�3;��tbPݐgX ��7:���d�ps=��4b���C|Od�N�.�gUz_C,�$\�^g&���I9���,f4NQ�d"����;�(gv�����fo:V�(C$�
���\�IGe�#�{�3 	�LC��RE3��8b<�՝1Ub�z�qV�������8r8�f9��}�_n4,�L4������pu=y�N�B�º�\eOJn��o��v�|�u.?�;�ﮞY�k][��4�"P��������Rm>ޮ�(@����� !�X ��b��l�3��l�e�~C$�Yd�}2ŎR��њ�(:l��Q�O:Թ�DH!��R�X:��HF�3��A�Yf�����1'�Edn�E^�>����8�1W�Ӛ_�m;��0��P7�q��/@uL{+K�Oc_w�O�؈���9���e���U~���X^P������tQ���^�{�
�(�xT�KAS>}ᴥ�3�,T��6��F�a�'�\�+��e@�h��_�����<�������nL4�T�4Spջ���ڬ��rk���K�Ɵ`W�1$�	j%����a�w->�S���^ߎ�->\���G%T٫�s���B�� h��;��a��"�W�>9R��/t��Ts�&T��at�ߞ���a���6�zCc��h0�݊70���%ָ�g�C�0q�w��9��i#=��k@�:ceD�����5c
�P!J~�Y��^f�K��ܪ ~�rC�����"чSM*�	�N�JFG�]jb��mea^����j8F%u~�����EWMӿ*ٓ�Um+$�G?,�<���.���C�{xg��j�O�|��D,,�.��	��k܋��$h�+�ȇ�M�'�i�y���1j�GV�i{��?��5�rt8�39Y���qӒF��ߢ���:Isd8�I-��3����}�PQG�Lȩ��\��*�^b �ē	����ݶ����*&��2�<�(���X�3�-J��lR���YFl��
��ˣS���[D��-��F��p{���̖����.���(���'�V�~�2Zڷ�ML���ӛ������3�gQ�� M��\>)k��G6���"~'%���Q�)���?���L�/5v۷si���(�b����y��V��R��)������P�N���ؓ����$^����5qG��e#���V�2��&��T'K����.{��K�T�d�1u��}��ca-_Z�5�]��JH�t�A���� �H�K?�3�쏫~I䎊�)���|�_���6��W�F&e��M�P.��j	��I�\�U��5�Rү�k�"�a��;5���	�����J��MK�4�|3r= Z�PH����I���5x$����SU����bi����#]z8nos�6�V�Wa�