��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ`T�}�w7�ɴ��劂�]���io�k?z��"l���Y��`~}5�LWF�Jǃi�wneE����E�j�2��v^��,��"t������s�%�R�����H�Ӆ�N*>\�k���dj���y���z��x�GS:�D�����QzV��W�2��%}�p���)���S�W��e�bd�<���A��{�������?�G~�����4�q`�U�V|9]�ZI�~����K����+T�3yO?��Wǵ��>+�>��z�%ƛ-��I*p�dc[�aI��]�~����΋�W�C8�-q���$�\r[�j'D��F��~P�te<��BKֈ;	j����x5I���P�a�g�������'+�AU�ּڞ�JbN�鉋��^#��VC�Ƚk�
�ҩ��ȋ�>�:ʎT������d�CK������5:BeUw0p����B�X��!1H1�����H�����a��F\��iި���w( m+�^c�O�������<ΓU�}�:��ű�鑽��}�j�b��/����;���u�ſ��FSH�N�9�9���]�?��5G�\�Z-�P=�#���%p�4���y] Ppb��y�4��*҂b�'PNr��ՈX��8�@@���mm�
�5"�!��Ҿ���Wʵ"^�FH�仈��i����Q��2!��5C��R!�
^jQ���s[���;	|��9�!)=\����]��_L�h�.�]l��ǗI8Xg`'~�9:B1�V'�b�p�N�B��-���ig�8`�d��Y��g�=#̲�>/���2���-��_����7�S�������k�-�6 \��!D���}N�Mjӟ9�a�ox��������8
�}�m�)O�r����by��='D��R�ਐ�V��3#���� ���'����&2������GJ��q	@�,-�A1؅%���HŃ��+�.`?���[uÌ�<B�M����"6u��wM���/ha�Yd?���)XV�#a��.���R;��M>u��mم���2BD�p��#{��[O?��a>������0�V��Q��8o����4�*iò��]���:6��{�A���:"�9��I�ų�1y,0�tǍJF��0��G���\��u����|}�ԛ����`il_�K���߳�倐L��yL�0e��N����n��������βK�5z ���Z����%�c\��E%KrQ�Ͼ>�&�R�H���lu�|�`�w9!b�#������ �>���Bm��6q��e �^�c>�~P~�Vt�:�҆�\��0�2�Mf��5@0�>�Y"��j�7��:�V��ڹ�Q�ݩR�q�ts��-�?��B�x��b���'@Z�e,ۇN�;�n�Ҟ�s��>c�	m.�����?�K�|�a���*���Vm���+)rP_P�%�yWˆ�$�@f��9 �D�q~�P]&�ҁ w!��G�L�٫��r�l�h�n}?�dJ�q�$��6�VM���K}^��Sb�HVHp��R��^�p��� �Ɂ�~D2J�p7��1l�����%z��}�����O���s�j��b��11�#���ϣ�֡��Mğ�_V|qq���m��j���r�iz�b�7���,�}u���2�՗o�[�v�u�GEgc0�$fq�@���g���� �:&{J�d1O�!<��V��}>�>�Ȓ�}x�"A���0n�ؤ�����ߦ��i���9�SdtË�;��W:��op\�_o�/K<�I+@��T|�
0�q2�Vgc�k�H��()�UH���IA4葳#�� �����O��� P6�D�B }u!�bx�՟�_k���.;bѶ�fq���.ehE_���<��|ܚ����n�<܉� ��C6ױ��|k2��)a�D�:"'Z��I,�D��)�El�#Ȉ���r9�9�d-��U��{M^+=�A+��ic�h��2"�JG�5�0DN��ִ�,���`���k֚������UC��[���Nս��9"NG�9hX�����V������
��Ŏb ��w#�_q�ةt%R��&��F@��.�b#7���g�����.�,�qoV-�z��2]j�K�$����Q���~]Ӭ<ٰR	;�
�"?�8��}��v�4�\�I�l<�uu���j��ևU���4���,�2�fr{?qނ-�#��2��dw�i�9$7�.��SƼ����E7v��D-���L()�Ȕ� �����
-M���K���C݉�$�vD�֦�F���ݏVJ�_�Z
�4�XT�T��D�=�
�r>�8���.�a���p�?W*�VB����quz�U���z���^��f�7��W�����+��L.��Q��`�-�0+tV��ӈmX��V��O��ow`ى `*C�ǡKf�Ɇ�J�1�%�W�6{��5�g����t���)���o���T�rܷ$���S���Vj3મ8+B�՟fS�i�k*n��I�t�	soX�Xa�"�W܏�wdī?n��&���Nm7{��A8�(u�����c��f�����]��K���'6���!T%�I<8�"�D*�s�
�u��!�BQF�g۞M�U��7Z���\lO���,#B�	�y�1o���ΰN�X��iN�G[��8��%̷Kd@�y�����*7*����R޼�~�h5�2�m�1��A�HF����0�u��#)��Ӎ�
r���=$��(V�?�,�I)���7���3�'6�X�l�ꗽۨi�3 �%<x�!���z$��4�t�h�F�Qst����E[��5����.n�p�>��l*�kdt��ә���le)yk:?ԁ�l�(���B��@+�K;�j��1Y�z0Z���=k�tw��D_,x��+]B�i:q�&)9�FI"K>�l������;�25�=q�Ov\���z�|i ���>��qTZj� ���_�@VB�"�&���Vs�����~�]QE�7�,������y��V���0�@��l���B�Lʔ� R^�ն@LO��=
��)�u��ԱX��bQ��?��������lnA��L1��lt�dn`.R�w�P��~2>�BHcE���1�H�+�~���z4-���c��6E��^� �[��g\+7a�_���x�6[0�Mmp�%�|+W���������P�xz����(k�+��bB�G��x�)!�T���tRfn���7<��"f��%�"o�1�Q$V�ۄעl��)d������&�% 2�8��d/�(*"=���B��5MP�G#^��͌��J�s�S^I��"m�����K��t�]��{a���J���`�����hm/��"~W�(b�����m�H�%f	?ˆt�h�B%Qm@������"�wV6%y�3���ӟz q�0�1���+�#%H� �&��ͮ�#��L�������0�����������W�ͺe���T$�С;�K���O�E�a�!&��>Ő��:�����l5��L�F0������H�����F���9d��&��F�_�*�[��~�"�#�����\ �� �u� ��*L~��??��p�}��� �)�T�������+���d���u㪋�X6Nm�GX��������GBC��7#�)�y�� �XD?���B�z���x+�P�x�b�J ��Fe�!k�c�z����b
F�R�uկ	r<k�ieqti��~���p�� bV��-�s���8�ߺ</k���]�Rf#gW`� �<A6�����_\�x"h�����Tu!:]f�R˳X�<@�5����m2Z4d,����wz�c�2~��(n�I嫛o� #�x�[�㍁N���|��.�&�h�I]���ب{+r��:����}�Ƈ��B�J��j�OT�-�t��2��<��~2X166�������T�kNvR���lǞ�Rf�3q����pVA�ā��_Nwp�I��.�j�z�S�X5���^�6����� ��@#*J\�㱡���ܸ랛n¼���W�}�D��bW���zr��YǴyZ,�u�Y�o�\����"Z��ذ4(^���(3��_CN��8,�K����+��JGt�,��lQ�@��L�^x�+�~��83T����M�'}q�5���}�J�p�kC�ь�nS�U�:x�aT�Q��SBӄ({�y%���2�� of���}�*L@�jn��h��E ��_ā�f}0
?P�IG:ܑ�XZX������?`��JzR��F�'�����縫����݈�!��Z+�`���MM�+����9�c LF�A�����Z1
Rv�N��Lh�h���&��1YD0������c!�Xp��¯(������L$���S���*�B9��6�I&�q�t��
i�q�tm��P`�ڠ~m_hN��1���.C��&E��1�0{��<��>�ֈ�ǹ~�dL)��b{NbK�k9�fj5�_��F�=��������^it�q��j���W��n��G�jO�%c>վژ����C6EWiK�y]�����!8�l����f��b���(��1M��w;�s�����εV�`@1L�fa�ti�D�2�Ѹ�(��l<(/=Zߵc�Ϙ�``��0�VcS�K,D����z�N�p�TR�?&˹O�nEa(�+H�1	�g����M<-8`�J|��M�f���{�����Q��5�9�Zہ>����9�r�� 1���X����r���ߠ�Ry�Zc�m��1�)�s{| �U��)�z���=���%2k���y����qKaߑ�N�4�MY*9�<z��x�³'+j��t�D)c�F���U�Pj��1��K<�c�6Eì���VZ	�9��Fޏ]o]H�fl�e�,*ak@V���P{T��e���$���l%�� T����#�E��5B�_C�8��s���V��6�� �}[�[�ǹ�0�9bS�G�~�fQ�����al�6N�}1�*����Y᭤x�9[&ہo��vm��W���%�
��B`q+�����AV���u�	V9��W�O~��S�zn]�P�"t����r��V��~_M��U��x������7;�Ɗ2Ľ
k�,"k�a2�"�Pܘ>M��>=�7�T���;���?�g{���x����w@�`�1)Ouh�B_e各t�*;�T����X�&X��8�i0��}v&�>�����;2�D���O�c��[�ʌ��H�C��,��v��F#Is�H���ߨu��� v�OE~0�)k�+��e��v����x�	^)?����CB?K5^(���:��%O���q�c��x�zT(g��X0X���[�1�p�Q�Ƈe���<KA���� NW3�ʔ%�|օ�c%�^������{���+�X��j��C�2d�#f �k�`A�h��`�!t��<���P��:!x٢ww���#���t5���,��X ��D���/x�BE��x�����â�L�#��7��Jn�T:�����rh0�o?6+���������H���ʼ����3)��M祷}��6�U�	}����O��f������[��M]����p�\���rM)�i�h�\F���k�c��
T:�X2�����BboxS<S�n����*DN�R�1��E���ÊC��,��>�蛹��H������ܻ��-؛\�CpvߞL�����jʿ��,�)�K�T*����q�d�	���0�F�l�]n �fk;�,k����sC�����л��[�f��@�n �(���1��-����R�Ohf��\D�mP��q�ل6<aZ�R\[������s�^:q1g���T�!��O`�"�?6� D���kT]�|��v Uv�r�\�NV5�;MKUs��|�ܿQ{��h}%d3?޾��Pis��Q�;��Vk����xd`c����88��t���I6��P�"kǥ����vm߅���-�Z����]
���{A�l
*���c�4�?J�d��1��a�u��K�vЃ�~Q=�1bp�˸�6��� �bH��D�^���1!w�%2��K��p41P=A��R�4F'Ҍ=;(e�l�G��}02}�G�ǂ�!Efh��(�"�r~�?�Y��H�a�daC|t�;\Q\�HT��
}t2L�Q2���mk��|��!3[��ݳ(�QWO�i��Q���a.��@�tXQ��q�V4\��P6ü���U��o�RÙ/��?���Fu���"U_[��)��Þ���])K;��{����kն%�����Ʌ�W,�x��]q�q��L-���*��`a����`It<)&.�Ml�2�7��,��ǈ:fa)I�jl�}��Q��䀹����
oL]�R1��3��k�ӹ�����Q���.�V���a��2A_69�/��&�p���%��O@&�2>�R�:�>,���yCsg#�W��2��|�5ۤ=�5�H0 �ҔЈ��q
u3������
�|��w �\��)�L��u@�R'�c�F���J\#�!B*�,��6&AU���wOB�4/��u�L�|y�U��nO��XD:�L��Z?U�K%o��5G��:^��^5��i�ԣ���,~����E�^@v����q&t�����23�|_L��"\��fE1�4Jo�O!h�Y�I^IT"s��z�j�� �D/����AY�hE���o�������Ӡ�,)��X�+�'L:�^
�z �4v!���^�y�3��|��)B�b�N1�)R��`���*�T��%����i�A��Is��v"��񘵑�s�}E��+sɗ�k�[yf���%?'Nxt�m���
��%�_�����Ra!���̹BFa$�%ΈgrV���T���_d��Ӱ^�hp�T�`�Og��%N�������v�K@�_�&�E�A5x�k�0q�@U�Xq4GB)'���d�~D��2G��벢(|�[�.G�h��g���S��%dg$�ՠ��m�#�����zR���e�4���>=��,��ҝܰ!dZ�?�}��v�eUEj�/��p��`D�>�� �sg��J�jvez�����dE��=�A�N�Ӗvm�����ǂ?�bvcz�2�"]�adC�H��dt���.2�����) ��f��<�4���9���68�IC�U�;C�Ï���i�J,���N�A��2(l�VC�<?7:��G�l���.�<%���t�n�
LJ�=�Q�Vm@Q��n�Pr��3�d�ٖ��JQ�VBG��j�x��:[1����X���	��3#����{k��k�
��'������zn!�laK��{
L��m�������	���,�y�����s(�S���Y�����՜���<K�g���f�qc���G�R.M��6�e����3�>�����/`"���G���6�'����Ew��<�RF�_�m D�� ��Õ�ط[���uU*�� e���-�� �0~�^��X�����Dq��?��#��������3e�B���BG8��e�ĸ�g �?�K|*`�Ή\�� ��sP�@ҸY�'.��~����V����a��/����v|p4��C��,�`���!_
y�J��Tܼ��:���YŠc��5��W�f/'"���P�%�S�Y�47Jw߶�DI�q'��I�<m+f4���G�`�����#i�<-xGgAƢ�ɫ�%"�`��Sj��qs�Gc��vXu �޹�'2c�~-1������2i3��i瑊l7�:�=)@�Q���ޮ��-�T�8���7Վon6B�8"s�,I뱖��5%ź��Vnu�	3-ew��>#{G���҂�^�t�}�3a��@}(��Ɗ(����2�A�Pn����n��Vd���_�c�����Y[�Pd���*���j�����mc��՛��V��yG4���D6$����k$���9�`Ͼ+֑hS��!�E"7*� !���7B��*�zk�qz���#*�U80�ɍì���(0���&��P����īk+��`\��2���F��&X>��"��� �݌B���#Ǝ_`T�@ Z�a���:����Y�Δdol��P��d-%&��آ�����X�;N��gA����gc�ѓ��� 
X��.0H���2��V�zD�|��|��,�Yv�f2�U�qۑ0̋�{f���H}@"oL�a�i�Ke3�Tr�P��
:ZT���{�^<8T�*��nj�@l-�:5�'}����8c�X�ฦ�^#.[N�8�Fg�ft)�^�����_�U�`��-˟x��<���z�0&+�����5�r�H?������2�����m�%Rb�;�HD[��2n��W��:A�J�y|U�0�����?��sR�xC���O�qʰ��R��;�E�;x��-	`��5��?(��$�fE�D%��ݜ�8,�S5
�9ޜ��m6�((UR����z���!�d7�Ph�`n
�3)�m�J�L��]�婁�p�#PW~g.f��̴�U����7.��	~�X��aYF$b|W��0�j�=��[?��T�t&.�¸�'"��h��S�3�'��a���.5��~��'X����:�8�X]K!�gJ��m���. �G7>��;f&Up���) f�nN�u��f��>Q9�+��Ӛ���(t��Uӵ� �:*^i}=�⑐�b���C�����4߿�������nBY���%�5����/�W>�r�T�|��aT��4Ta+c�?��������OD��Й[�:�.EU��=��5)Ԡ������?��);�Ӏ��d�Tl��g�
O�z�)�d�VA[/t �H�5�Ŕ���%���xT��XT8@Pn�� ���ͼ,�!���U���R7��89
O��P����nó�6F7����,���VT��R4-����� �E�Nk����V�g� ���A�SEkIҝk�&2�$G@6�;}�F"��+�!�%�b�_���En�^��*��f�׈{}B�ޒ�����P�O/]jB�Ph�TL`���i�a��V��(�[ѯ���O$�.�n�f�Ӱ�ҥ�oJW$��a<��ĽQ���Ie��K��<����l,"��4^z��h(f��q��v���]�0Q�K�� �̄�I���ڼ`��i�f�l*HotO�#��ܭ����- �<��c���2�M�$�
��dͨ�i��2`�ğ�-I����G����P�̧8 �>��Y+��kQ#Y� �Iԁ��R���y*��}����`=�������es���KU�`/�V=�p�X�c<���ֻ�EɥP>���Bj6���4�P�-'{�[Ct�`B�Ez�� f9�����߂�u�\�%�]%��<,*�Nevd ���������ۅ��L��_�^���r��P$�%lM��	~�-K�셃���a\���}y�)�X���]�s��3���� �t�)�OD��ɰѭ�` i^9���+�ʦ�.3z���%� �.v��Vb��a�L8~�=��݃{��',p?*?�$��z3���s�����JԪ���^5fF��MO#;�V�Pd������J4P�(����l��3{��L+�q�lW����� d�!�<5��J�/F�'?��S!������&��*ǰ�A�K��j`��@�K����)ָ8�r����C$]�Bc��yWGq�� (������R޸S275*����F�HC�ܮE$[W��_�*`)f�d<��2/3��3o4�2D��
�x�z蜹�'�ǿ��	�z���Td����bV��`xHW�Sllq��c*�D���sD; :ڿ��(CSc}��sN��i-�t�,+�a��j�*3����'Y�P�t�j-;���0��DI�D�1�Ҩ���S�̈́���ҕ�Mm�⯭ƆD&�&�Z]}+�]Dop���"������'>�ً���]��<NT��&3��c?� l�zG�@Mk�į�n�$���}�8�=eQ�( �����I|�҈�s2=�bqDzU�|L�![�H���p��s=ΑHR o�U���>�+����[}=�	+�<�������T�w��*Z�0,� !�`y�6IΐV�w���#�H�H�S�����&�B��}~�TN�Åre��&��7�/��z�Ja��/�>j�uǉ\i�����~��24���S$.�fb��!~�'�y(�����"&���%ы�9'����S}\�쪴N&?���8N9��ڣ_�[^bi_��j�c�?-�t�B�x�P��I����f�#�8��H-7��߲����V���@��U��W/���1p������VT6�����m&��{���3�.Wb���.�ܕ��X��Cc'qJ�R2YHU�@�	�f�ǩ�	��,]��8�8;��c+ۘ�K{1�i�.��4�Mt���<kx'�`�
6b6�+��"��X�Ltd$WY�	-�,�2ڤy����pݵ�$�<���1a�m�a�ߐ��p`e<HU�P�����,�P7*��E�+7
ɮU�^ Γ�e�Z��S��Ҙ8����c���[�Ueo_%Le���^pDS|P���Ĭ���I��/ L]��K?��<��_8Q���Ihr�5f:�ͪCiB)��`ء��@��g��.^�L5�T��ß�)vFy/Xk�혠Du��F�05"G�.ԅ��SLXc	B��驚�us���['A�w�]�@g���An��#G�e��u�;�٦����M^���DnY���aY�Tvە�uZϻK��>Sw`�:3i�Z�bG�p�x�8����\���q��W��Z��|3��t$��IN��Ϣ_��$�䬓��Rp��v�Mg�屯m>Y9��[�eo�`�nQ�H|q*"��q��ut���ԬO�1�6�����_���."vg�l�Է������ޘTk��K����9���S���vɓHr����S��^0j⢬a]j�M�SB>I���S��]i�C�͕n�{ugϐ�/>1�s�ʱ�T��C��T�= ~�=%)R�7q��R���h`��^�*4Zf������z��5rd�〯è�Vso���C��͌���1�7P|���/��ƃ�lcA�ն�16�w-ӵ���AWGW����Mq�|����c4�t��*j��c,��o?q2Ʃ?���>�p����7"qT|`��}��+84{&fr�ҋ�Jz�m�� �xj.���|X6N�>�h�nX ����#�
�i�6��uH�QX����>��Yn&�����@V��PB�8�꣢�4��g�m��:����5B慫iQ��Ϛ	�$T[B��TEO�6�&���68:?p$��ɚň"�yw�Rb$��'��(c�p?��O�ب(C�<k���5��DH��MU&�F�c4�����5Zb¤,��G����z�߂�E��,*HG�i�UkuU���&yv�|�?!\׏�w�FŬ�{��E����������ڄi�W��
p��'���E'���~S��1�,����\i�ip>�#��x-�b�y�Y�p��׀����E<�$}5E�.���}��I%.�[0�:L!E��Q�$� Ǫ���ɧ�zO�ӣ���X3��g$����3���)&������g�;rm u����۽��T�ޙ���A� �r��8���|�OUz*��D�]<묈��S�<��ut	�r���e��)M���O�+�1!?&�c��}_�#7���"��	I|����O��Z�᪤��±��g����t�?���Vf���#� =X��&�$�W��	���=�Հ��54b�晫%z��ϴ���f� ؂)]엿U��*����6
pe�5'%ƾ~� ��X�^��;==�i-����>j/�עW&:���|�C�G�z��<1=��RM�����]�W}S]��p��z�Zݒ�b+b�z�c��
�'L��7<��]&��i��~��73�2��F���5R^%@���vm�J��%S.���.�B�1�=�X��%��=��X��G�K�`t"ܷ��@�e��b﶐~�c���ӳ���)W�@�Մp� �v�.����\7�G���֋��fK�Au�n�[[������̌x-U�P���I�K�,�z�\�4@��#�$��#�[H׏�W��?$쭚�I\�蟐I��p����%'W��R���Ȅ�މ�$E4����E2wZ;Ύ����@���u�4�թ�ߠ�倈c��|fψ��� Ь0X����:7��WP
u'�X�9p|{�!t�����%�ߗO�9�AQb�>��
9z������VG��6i7����������y���wz����a�>Zf��	\"�I�\��05�FZ#KC%i���"��=�!�A�t�3��0����a@M��
���S��^�P�}��
�b����Z��k�kH��e��M����U���O�ح��H�l�d(qv��Sj��N��K^ض���tz7/6��Pզ��?	 W��t�����?�,t.��I����7n�n"$���P��o: ����&�Ǻ/�~#���J�1ɮ�ǃ�,�����`
x�߇�6V+�a��#�\"�~��\S�¤�2)��S�`_���p����n�� .�M��ے�.mze�$��_���8���[@��X�2NWd'�Dv�fME�^5k��`�/�2e]��q�5dѺ#,{rSu�-3�V%��_1�8���5B�֟Q*ՙ��Ǟ��k?�\�&�Y�_J.�,m�dx��Ugޣ�kG�y���:�%襠K^O��eyw���΀��@�-A��I�Z���e=�yG{#�>���Wb�Ec#�<>�`h��P���u���R��.����]k!�e�<�<P���"��9��X�Y��F�o���	lG������� {yN��fz��_�0�Ԭx�d�%⅚��t��xr�B�D���/�U�0FK�s��$���6�Ie�jhCo���}� ������m|������HJ�g��,f�ۛP�GI�}�&"�/����n)�s����*ގh��~aY�Đ��o�D�UD�(�W���o�U*d�+s��O�β1�O�ۄ�S$�Z9g���j��i����~��À�'Wo-jvd�q�Z|�|�֊���S���¼��9˜<j���R��Wo�T�׻�I_l�oW���&ri�LM6�Ý�:}��s��n��3���Kʜ�]�	�B�O�ӌfp�<���P&��Z�l���ѷ��La�Κ�y)<I�o��u��Aa���&�8�i��䒥���K3ܥ/sM�e��$�g��@�6�~��hN	^��װ�����V��k0�H�w���V0_�K(L)+)?�?�9V���V��i𻌢i���> I�
_l�F���Jn����P��`W���Ui���
Ɉ�8�|I6�Z�(����9��=��E�C�E���3�\��2�e4��}]�2��f$f_���l�II���"q����g}ض*�����DG���U֫��!��.��`�փ]���|*��Gl���^5�}4�j���>�VH�V����i��SOp��Sʱ~�.3,xu�>��K�*������b��67�Ӆ 8Kq�Ѫ'��|����qHx� /�]6t�Kh��EFJ%5b����YQ7т	Z���+�kX�m5m�.欶%�~�I��h�@�9��k���Jg��񏶴�	
>�� *�S���KI�<�4�����?�I/9���[=�o
�"d�̡��
����r֡�x,t��IP�> �]¤��F��ퟖ]�C���̢�7�����K2[�F;��L#�U�i&��7�^�w���t仙�H5����UoBf�[�o�5<0kh?���#�HV�g�G.��&Nq2��Ir�pcÀo�3�a2z��7N*��*��jg������t�fV(�?�#���H����{}VogJ�fDW����!�8� �1�
�,tl���0 =�aS"�k�Eϐؤ�]�������,�����@S�Z�	�&q_�'�ƕ\���l{��EhC�V�}?1�y��dX㰺*b~�!h�i�@sAr׈���E�M
��I>sN�M���J�4k����H����HG�󟥄"�4��?Y�D!|s��*ik$
9J�9⟄/8k�b�GY�Q~e�	�sl�ҵ�L ��	i�"���$+��@�m�TF���1j��z����iV�	Ӆ��8*�!䊺Z���X/�m��k1� �hqe
���+
 #[��JHH8 >z#�e,�x{V_��hɽ�^�zYB�;6�#�닅?�Zi2
�(k��l�;�U}�����A0�J�0���vq|����XG�p��Bkj�{�`T�\��GU#��!a��*�H�U����_%��N\y�X��q0�m*h�v�ۤ���L�l��}���:���y�C�[����i�Bg�9Ց��F��_zm|�� �o[���Ѓ/��<��wA�e�[OYd+M�;,:��Ό׸ ��W0�������_�]�W�%A�6�\U��A����Mߦ-o��ťJ�c��{���57�~�>|R�"�Q7bo���hm��D�4�G���;�wB��<��I�?��
HB�bW��_��l��y�����[t��*J�G���e�8A��$�@�m�����eϓ�,�Il�r�Z�9��	�\��W�(�NBm�N�N���c����D�u�Uڣt�B�ll:d�	P�v	P�a��{�&���.�����z>)�I5�+0�� ���,H�jԣ�Y��&O��XI����%��֡����ί�,_�&��'~V�`GL۟��ŇJ�`�z�Ⓑ9Q�5�Y)b��?U��n�
�[�9��p0-��y��>�jUO[Tbh�'Y12c�>���9:F�D=mR�ӎ�R"�� ��k�����t�$-�Fy$7y��@7d[QG�R�"杠#�Q<��T-E�SX9���$(�e<f]B	�"��g>.�����dF�:�� t�5�^�V��`���H�Q`��	�Ak1NZ��&�ޮ�k�0��:��$J�w����3�c��<�"?�����PJ�e�b��G�<.�ZbCI>��"?���m�"�.���� ���r�]A�����k=�eye����)�ԡ?*�͛X==�������K;��W"��k�&�<e�X�y^,�:�aT�	��GUZ������0&�������AF����M�U�=^#�9z�x��-o2�,taQ+��T��LP�T���|xnT(���;3�CE8�,�^�>I�����\��@((9ÞE�s]�>c�y:M�'��۟c(~�
P�:����7���d*�ф�2�����ގ� %�;���S2���7�y�%�Ӝ�:�S��w(���ݼa� jJ2Ν�ĜSݒ#X�\	������8��v���u�����`4;n����}�̬�b�K^m�}>w��aX�+C~J�v��λ��TqS�R터>28츁~Y,Y�S�,c(%���;�
̈́5'-�D��ΌH+ѝD5����qeĽa|�>�w�#��x^m]�r�o����4UX�um������&b��/jm*�\�o��v)C�q��������K��ע�����G�\���7>ߦ�$`CY�2bN�;͘�5��׾���u$�e�U�z��X�{��>҆�,�7��/�:##fE�⾌�h�'MVe�F�!T ��Bv\{$����`�<�7*�g��%GŮ��ږ.IT�.H�Ed����	��X�Q%�D�S'{�a�G�b�X�h�V�Z���9�����u����ӿB�d�]�t�&�m���eǁ���qLo�l[>ڌ���®��JB<y6��0�6���C�o扞��+����\��1��k K�J+����0M���[��s��<�k,D�_{�A�(��;��?+��3���MA��7��O�i�X�WA|kW�Vp�AGs�����5�i�Y �a΂�<�V�T!^�V�j���нXV� � ���r�;��%�Ȭ[�T��[��}usł����y�=s��q@�e���<`@�s/�[5U+8擌��>?rxF�j���1��/��KS����ʤ�s��&Wt���a�4vL�vq��������ǜ͂����t��y�5�t� �*oPa�u�
{)���/���\�|ӎ���|�9�*-�������I�<?�(�Q�	,$�M��D� Ç6񫀯q��2�9+W�"�2XӖyڎ����H��^I�}�:�t6CX򑮄J�i�����cmv���UZ�/��v\95�9��3%G�W����M"BU��A�@�k�R
ncH�F���*1$g"ʉ��%@]	F֤q��Ÿ́K�u��G@CEM�B��&��R/D���7��uX�4V"!^��x�7&��1�$�L2�sܒ���,���&�?fw{0���/�~��H2�xZ��!ؑޖB�oC7�11��y���~Z�}��e�~��6�ɨ�GhG��v�Z$sk�W�BC�E���R�5��OD�v<]E�g� ��y�dy�jK	�)Q~a��Hk1g��x�	��P*�z��U�s��l����r6L�������!-�]rq�K+A��'Mu"��?�m�PY��I쭀�d�����E}�(_aV%�������R\���l{H�����A[�E;{��⺶�*K=�굪|5�����Z���>a;d?f�O~�E�����Z;������@�e���@VP�qQlT��r��A���۩w�-a0M�y*�J+ ���E�H��툘�F ����ı�W@x@�v��Yhs��<��V���X3GyU������N�X�����~u�\ T�F�5�Iݜ6��>�{<����8�'Y�^���KL��޳U����a�=��ݡJj{�`Ud�q���kJr�[}�}��O��v(ȹ��34H	�kP�	x��Bnb��)|鍶����R�hY뼼�#.-akM�	L��(� �dUG^��n���"v@�va�.FY�/,l���m�\&��`hdj�B�'�X.��@il��/3hl��9'<͸���Wv��{<_��^�
��
��CkUϞ�&9i<S��S�+��m��k��j�%�3}MF�]��F>] <�"��"p�Cq�8�߼OP���1g�Փ04���V��E%p���_6��Fk׿���b�ZF��z>?�	˯8�A�e�ލ��#Z�U�b) �ه���|'J@ie4�c�����-�K@����dgp]���_�.]��E(9���W�
O!�[܌G�F\97����!��$�����!�)I����klm�r��r
�9I��+��&��>ٮ���C�fD�%��֔C���Ql���A�R�C�h8L�X0��n��D(�T�]&�q���OA	����ɒ Hق�F�xrX��:���8���,��HH��i1r�e*�xϥ��-{�E|א�������.9<0��d�$pC��?kÉ��	�-�_�fIY�h���-����b�s�F�w��U{���)~����: �nZS�T��+�	���N\��X>y=�n´5�_lP5�Z�˙����J��8�K�<�`�/��Y>��'D��>ΰ���؁;?�xKC��E'��ū�A�gq�����I,i�	̈לp��hm�Ԕ�L)i�cG� vTA&�6d�j:�����;��^oZ�ktTg\�x���ڑh �L��~,���m��LY��"nXM{�l|��������c�(]J��z�i7��Dlj2��1:T�ey��ch��s��&�Ěe��R�����5���^��_#���SnV��%����} ���x>h�/y��=2�"��������1�� /m�A���ﻋ�CZ��y��l�AL�q(��e�!�Z��80��j���?s@�gL{�s�7yvҹ�.�"�ޟz��M'̴���Tr���U�ੁV=Kk��,]߽G�Kr,�a��7�ˢ$��\oۯ�ݧ��A��������ʝC'�D�S���Z�S��!4fV#[`QT랩���'�L�N�)/�h�al��:�괥�+@o��裦i9Q�s�n���F�B����;Ç�}��ߦf�E�z��u'?l���Iy6g�]�S~���Ǖ��X��K��l��7�9T\�����J��7���vOb��5r�w��l���W�͡����D
��w�Y�#4�B�BF �.*�D��< ���+B����g���Q�a�DvІ~����)'��A�0ݧG�:���ϕ/H4]�)7J�N��7�	�����ބ��o�E���2[]؞aD~d�� e�&��AaG�JD��o�X���ahKxgƤ�X'q�F�PL�l��,�,hK;�Uس	Q!ݼ����#��n���yh��~��S�Pk_g���[�d�Sj�k�0m}��3|?}Bf=�O?�W򧎦����<8�C�ggN��*�6y�j�����K���Q��x<��z:��~0��G�~F��x�o���P�R��E��ܺI�!�/õ>�zHÈW��ۈ�P��"��>�S��*��Q��x!�������� ˄n`�\����4mL��Q��	O�>d/P�?xW�H�+e��#�-�I�_d�g�Z2m&�d��8�Љ�����/��O��ٛ?�����Z���&�Q���A`�m3#�B-LD��n���!o� %���B�6�:���򹳫�ƟJ�%�+B���xQ�Q#�V�׌�[���%WܰsIhp'�'�ц�X��8�3����ҫ� ��|�"�L����t��j���ӯ;���<���o(��x�7�_?�gi�+�>��p%�nr��e���SM��h��J��}��>��Y��½��9�d��v�"sǬ-�O7�����ܲwgwg�`������F�U�-����>'r��۔U^��8(�, ��ArE��H̓�9�;�x�az��~�aډTvceq�=���S�	�Ď����(~(�Y�������:�sx��ɺ��f���2�eL@c�w,]~>!44���u�Z������;4^�Z���ڪ�7^�Mܛ�l�ï�QLdT��� A����b��J�/�u!?"�h�.�����W�mR�u�U>rj��'%`R4g0) ��hr��¶'�d��t��b-הw���SJ0� ��p��h��K\5�����ۓUN�|~4��j~wp��Iˊd_>z� 0�⭷/�q�JA��F@9����x���xCWĽ!s���s��V* `����o�5@)��EY��۷���l�!-���B~��b����'m��c��(�_lo�oGK�^3;���?���kpM<4�<׏��N��OD���=7���� ��'��e1�eN.Z^��0a ,��W��JE�z��H0_d�?Q=�~��	xtۜg{���A��/]u�M�V��T��R�	�dĔ����`�Hi�+�e�p�n���������U�lp9n����l�=�9f����"e���:>����ܜF������Ң?q���&IN�L�W�&B���ZH�24(@b�JC�P���� ?pe�ъ`�H1�%%�6���L�R��붂��6z1a�[�M��j[w[p�&�f�\�b@n����b$�ٝ%�3��W�������A��lޛ}~�WQq��sEO]f���p�T3���-q�q$�`�ۯ6�&U9l{�;���׌�����Jh�)�ϢxBa��/��7�ѻ���0�����д���h���]�l�,���q����n3w>.�%R��)���O�9 %�6���Ǟ����nN����2�]JJH�{�9��:�m���B���ΔF�̶j���B^���vZBGዓ9�����j� t�7�k�;n�"\M�(Dl͔�W��� �����݈)X.u�fX $~�IQŤ���})���)F�6��ߓ4��A�ECL�?>�\����kW|� � LwѨ_I���f/�I�@������1�p?��[���j��_�y�!��k�����֏y-��
��7���9rIwsl���R �K���m�UF8���#UG�ɥ&�]!fOǿ�^���yd%`�t�P�=)S�������Yn*iӶŦ.KI�=1��'}������uʶ1�&Y�h(U��D���3�*�>��4��T��?�֕�L�~3�gR��C]C�����'0�`�8%<�Sbs5�ܬ^-f�i'1¬j�o85�~�iR�k+�P߽������Q�k	�q���V�3��F�e��)���b4ˣ=�[��~ ����ֽӖ�n�?E8Q��@b.��3�����C��@A�<9���{�L^e�
�0~4�>��`{JWcWvM3_n�L��*�3�=ذ��H�~ʑ�
a_ˎ�f���V��6x�o3��[��)#<�Ѽ��+�[BA��|�4�e���W$�V���~��Znq+r��_�"v�'�C���ª/�c=�Q��4����U&L9��s��cE�|"ܜ�P��qc�%!�� ���`<W���ҰkFQ�y���Q<��EX����Gy=�1��+<[w�'�x�䖢ɂU8��B��s�-�"��Asl'a�E>OIB�*|��D落+xn�~�k��~K�5�m�O���W�}y�mk��-��b�<�ε��#�E�j�$Z��dYt��&�t�C_����U�����C�W��7�-��$aՍ
߫�>�=�3+�}r��p�t���U�3;��!�8=�h���v�a��������-|'C&z�3�j�:�YEϰ�Ady���6E;�t_A�9J��Y8�,��V�t\_��$
����C�7��9��^�����ˆ���<h�����K�Y>F?Ow�r��ܬ������"�J�7p:W|�����O���O��dq\�,r'Ȉ��04!�q��w��6���� V&�+|�p�ˎ2�2ƽ��)v�3d��7���ݹ"���Z!��ɟi�'�B����F�����nkj+S��TA�	`�D����!#�n�+��P�3�u��aA�r/��9ƹ��h�f�Zށ��&,�a()��B)rT#U ���'[�溰�a����7�����h"�t�uiB���Q��z�3��m+�5�m*�-Y��n��ю�*TOw��w)�|<+Цo��0��t�u�� �#��urM�L��2p�P�1D2z�3��(¥�
��;];J��+�tDm����3��F�A;�)H;g�P]S%�f��I}gڰ����A�/�Z\cV�e��SNk��S�GO�����/}�1 DJ���Iq�<�șy!3
���	�*I�D�Ɂ�r�cD��­�vX����ҋ���zn깝��>*����p'��A�M���E[���E
�#�nY6hZ��[��*�ZrDBb�BU/M��Fe2R#-���z=Oj ���� x:�hL˝��3+'b��-;y�!��F�˓U	�e��KM�K(����=�C_������y(�wV�n�[�Rx{Ѫ?Uf��un��1��aE�o�M��e�PU����r����~u��*��T
�2��_�RS�t]r&pg��/�idW9�>�<�K���N$�����aᩬS��X��{�6�H���·n���m���	ل)��e�]p5�ѝ<�dľ�1��|��WX�&���!vT���;K�>�e�֐"i-�}����PD\Y*¦�}��X�6��ۓ�ԉcc͏�+���8E9�����Úb�#�yc	ȶ�C0�-���p:�\C��
7�l�ra�?�Ꭳ�_�����8��>C�i�Pv�VK�.\$`����[����K�MXlev.g���s�xhQw��@�iߊ���:Z��s9�`��
��t�t|�X��!���� l^!���2�,8�"_�:ta���J�0��4+�o��t�ى��G���bË��U�mң������X���>J��z��HR�q���V�����V�vt�����4/#J�Y��]�sI3��،�(�<�dۦo��%��'W��[&���p�th���ҁ�Q��!���?���i�/[C������^�7p�-5Ih�����������/Ј�%4x���{N q��I�c��p�kh-����Oۧ�1�u�3�0�0��yw%b9��~i�����J���I�H�%u�$i����H�;%�WqM\�e��8y����;��I�Tw>GF��9�Gڼ�=���!��NaA����$���h�r��枻�I�Q�Ԙ�#�8Cá�@*s�]Nu^H���^���[���ƪ�b��X�"P�=�(����og�J���fE����x�|Jm����4C�<"X���}f���^.���-��RWA�P�+8�d�>��;�����$�b�<U���b`)UP��3��C�FK!u��*� |e��DA��=�D�����M�M��`�o�-ځ`�.�=�_-7t,�k�F�D����/��Z������4��s�xu�0�Tw4d�0��a�M4{xh�ޤ�
*��˃�M��@��4���Z��G3��+Z���O^6 $����}Jc׃'���L�t	��]�8�맩����7D�߉�-��l��TebK��F��0��^?��M|��.�$�j�*:q�.�Z����r��0�iqMK��p�+ʺS�0@���fzέf(�������3�/;��Ns�9ѹZ�/p�`����xi�찪��u�h�ğO�bfw��0Գ�d�^��-�C@��W�������(6��Y�%4�����_�{�W�>����=�5*@�H[��;����i�X�I��;~��[~�����'��L*Z���)���I������&-4K���\Ā�'�8Z)X�?�?ׂ��P�[
�rb�+��Z��4x#~�=e��_��y��T��&��ud��g9�;�x��Ugy���)$�F�,΍��ն��PE/��z����&�\�33V0�O�Vc��*r��#,����@Rc��	nu$�4;g-8���7�����|��	"RW�{l�pB��g`� /0愷�_��@��1��;rz���0^ѱt��`��U�̂hP\����A�W��!ۦr`�U���u~��*(������W0���zv��~e�$!�����yz(= �c4�-��Ĺ��r��"����JN���6eҰIe�P�d���PWZ�|4�ۡc@��3�8��k7�i��ߤ�U$	� ,S$�l�gIJ��T��)ڧ���c�6E$PGU'�7��lGYv�S%s��.����m���[�oDK��U�#�.�Pu9O�- =v�\'�졣�s���nQz��z�ó��0�JKi|����L����]�r⼍��H�߰����j�}=�X�B�dى�kT���ֱzܢMT<�Uk�8$:��t�}����xK�k�{ԡ0T��ݺT�@��Vo5���O�TD��l�N��!�p�{)i��6M�c�F�����������Β��Q�\����(���%�b����
&��M��:���g����Qw�м>%xJ��\t��ݠ&�}����Ñ�(�Ծ]��)ӑ_W���B��B+F{//3�u&C�Z1-)���e��:�[M(qq}[�m�	���=K��i�+5x�h;$^1�v��������+NxD�����4geE�r{�SGkoЫ�-e7�����L�F�{B�uO,��ݪ|�@cJ����?���r�*'p/-$��K	1�ղ��ݪS�du��y� N���Naڿ�1�=�2M�!���W�2�3����-������Iؖ�ϙ
����JA��@��\f�U�F\F�m�A�Ab���W����J{��E��L6��r�V=��[>�N]�h_)���Ua����������<�^�Z�Ou�o8��Ʉ�M9)se��~�ʁEʫ[��3�O��BO���݃��e�I��?g�N�����B����JDJӋ8å��n��r���j:��	,��%�Q�uK����6�#u�'��R�^��@{K\n1�;iPЀ�0�5?�����3ŕF�S_�h���ʒ�����d8�p�T�A-���M��n1�J�M�B�|�3\�=�VEk|]�#q�@��la��C�1�ws���$�ԺKJd�f«�/b�B�D������V{`�v��V,@\��G�aNm�ù_!7�a�p�Z��6��q�g"uj�G�� zW�и�J�B��8kZ� 3s�mU?(WW����0�7G�I�*](B���@��"r���֜�e���2�e7�l1�
���� fB�XolvP� �8��<���i�Ǻ�م��� ���~ m4Pv�^�*`d�QeDu4��G�>���z�h���[ EOUt|�>W_<�{`W�;��� y� �� &$�����RCT)!�;�L��8��R�r{�On�^�yTZ_�(�4'��.�ty�8�����S��C�H��P�O��!u�~��7���y��ߋ�Vh���4/䆠顫��A�*&�^қ�}������6=lqٯc[�g5o��KnHw̍��J�����|�ah (�����CB��M��#����oB�B�o��F�\��T�!!k�ďΫ������}%8F��)�0��{<��%�k�1���8�X#�njo�rCT!�&D����>;'$[.���7����G�~��i�����9���g��������"���+�=�|GS�u~�Mj��N.���f�]���;u�HX���R.���y�[�>��:!�W���L ���;͚i���?O���RDFi_m��jnoab\Rw��}��"���z)��E�i�ZYp5���2������C|�� ԭ���Q/s5�D�9ΏVCK�Kq�� �lB>3$i�A�T��A����y���z֜e�~��e���b���&�Z4�oݣ����(;{vj��&q��#�P�"bf=%6��؍ur����'���>����,R� �p�c����6�!`yZٍ�!�.�f��%�h���m|�<���|Y���6�\�ܪN~Npa%�����̲�����������ῂ��i�t?:Y��Kub�:~a7.`�ƈ�ZV�W�b)���|t=�|8=�K� j�$���V�nYT~�2s�m�|�>'8�kh�^U�ӌ߃~�Ss@\��;�n��	����rR�̬~���%̉H���� g���΍������;��m�;%C�rH�+;Q��Xy'"����<Z�������1*�˕�$(�K��/�?�R�DB�S0oN������J����d��:���;���G�r�m�J�(�Gq4凉�?�|$(�omP<���>�{�y�7���k��Ʒh��<�K�젽HD�K[����ց�^�TM.S�$^�V�8b&�G]���'�$D���hCļ�+���lr%�^� y��
5x�0e�}��UY2W�q� �}�E(�O��͇�,�	�ml:�
��m%n@�Ǟ��[�	á*B�(�����öL}�L!�Y���)�͑�J�f�ޫS��*��ϑ�
�yL�1)���H��^4|!y�[�X��ݷ�r�� >ID�t�*��8*�,���ߟ�������^l�#@d'�o>�b��_
��5���	��*#6�7�~�h��h�|⸿��݁�;�|.�A�p��q�,ee-��#fS�G�)D���Ͼ$h`i���_t�k:ga�������+0 �M�XR[A`� ��o�O���QjjmRq��✋����9 ���y����[~G9�R�af�Y>����uÝbŦ0����yy�?q��Q��Q�tB��.Jd_���+�PBL�xE<�d����� �T��B����/�(ê��x����<�����K2^9���"�j@�k#�����;<��o�d�L��E���ZT`�ƽŪ����*�3Ǧ���Q2�@wX�<v�F�D�a�x��3�Q"*g4��m�1&nbMk�o�>��0̇�I�~ ���Gx$6��,_�[.
�~pS(�ɒ�0�q�f% X]�?��炆���h���AR�6"���� 3Z�Oe��aԮR0�n���sj�=8*��;S$�ŉ ��zm��ʔb����ң��g4��䤁<Ʀ1�'�"x�1���v2|˷O/��!i�x���Ճ7)�$�f"ʺꇳ��?�iz��@˕����~��6���!#r5B0,yGg���I�U�� ���!D ld�t��t�]A�!�f�_p| HwX�"99��"��Kz�Z>�!���) e}��X��^EhO��������t�h.���۱�U� 㪫��U��>�F��$��U2b�w�/�	�]~�ҭp7��l�K��`�}[�h���C~jQ|�7���#���Rd���U#ݪfН9R� �	�������v���6�"�������E�/$U�k���K*��-�U��D�^�I�.%*e��_�u�����v��
*G}�u���n��=�����.���5*���L��O{j0x�XOη�1�WF� ����d�e��	�s���FH����
��kIJ͛ɫX�l��T� ���"� G��?�aW����T=s�O{ ��=�6�%���1Tp�P�4%�?��V@�ͳ�+^�����˶F���,0��xV/�W�A+����3Dk��nK�� �lҐ��o�G"����X�Pog���X�^5�DJ�����J��Щm��˦Np�jr�8o�K$�n�_�d�,i�ʎ���͎)����Ǉv���0H��  ��µ�\H��g|@����hP�G(݂�]|����ݬ�0���{��I��|�mY�>n/��@�\W{x�m��
��uK0������A�����u��l��Yn��Q�!;8]Y�%V���v�%�__?}S|~��]�����cJ�|�wq��֍#-��o�m?�Q�R�@��Y�d�J�j�ś5S&�]4�%6�N]��7?�
��39��lԝy���U>κ�r�q|x�6��k4�f���"B&h�D�wP"�f7r��c�"")B?�X ���0ݔ}�֠� :x����E����w���v)�c��L�D[�����H�	{3p,�ډF�.�!�;���P�ј��}����ƪ�0,�0Hm�|����?Kȭ���g�d޶#$��o��JG΃��A�$�9�l�d��D�H�������M����ۏ��d@��Z�c�t��s��	dƼ��A��m.��lT�6���u������Z��ծ�TN�����et�QD-۟�=��r���1���@����k����S�꽭!����H��=�arwu9�Z�%�SPh+�2��-�X�z!��c��pe��X]�9�_ xqi���-Q���N.�Mh�^ON.�ߓya]3 [JHٮ!tQj�"�w:'r�"��8~i�y7	iy�m��=�^���W�惼.�G�j�$a?�ߚk��T���ZvUݑ�%��d���ǹ�\^���܏M��j�GB&8d�?e�S+�����&Ak��"�ȞY�Twܢ�,!�W�MVm����2{jd��4v�/�wx��������=��L$a{RQ#�/�ç;:�wZ<O��X+Y�D�՜F)i�F5ιY|�a�釱iOu"(�9�nc�!�(�{�ZL���y�^&Q^9'ص� ;)KVp}IB������5���^ne�4�O'�^JNU,������J�*K�O֎XL��k/�a����	��R'��fذ��B󦮻z=A ��;�\�K�wܓE�\1����L��i]����F���P�$�*e��\mD�/�ӝ_�NN��'l/Y��&%P�kWN�e��`n�p�n���aem%���,-هn/�C��p����9���ȼ:i��\�z�[3Ɛ u�[��R���-X� �cR�j�=��K���u �p��=wVg��SmZY�N\:`'���;\hu=��fL	���)	�{�U�='� ����K `���p)Y[L�������T-`eL�I�0+���C�2(��5�W�{��,?��z�������e���o"��S�rW7m�,,�Z-��m/���
d�B�:5��@�
G�o|�^F�Kqe	��s8�Vq������%X�b0�xg�O4�3�۟�>j~�~m9��`D�?�oj����T���C�sw�Ԯh����R;�Q]r�wi���oϦf���IU�DKEq3t���lw�hX�?C.��6��7HD/�0f����-3������E�2�Nν��U^65�L�|S�����^��]ѥ�\���H,�:�U��Q�����?�0�n�+#�T%�:Ryg�(�)w�zM�`M�J�Z�<�v�;q�{"eN���&��[�ܝ�dE�ZZU�Ж��B���y!��������@���y��T��:��n�K����gQ%�h�n��S���|2V��'f]�����5�Ƹk����xg3F��ۇ�zػ�%��z��9����o����m�1,~F��[��eD֜Jjw��z�3 �y���Oc��;�t8Cid��uL�Z�z�%�U��IfEj�.Bn?,Q4���R�����tǳ]Nv!�G���"t��#MNL��0G���0(r��gJ�o���ZX�3�����M	�D�W���v�Q��+�Q$�!�?�B����]�������A��Q�e�e�N.L8�t�D�9󂱴n�H��e���r�/��!��D����n��{��P�j��
�������>#iۘ�#�i�#-kE�	m���Ҫk/�>�����\	�f ��1DS�:�W
L�Xf�̈2�jzCdQ}Y<7��/��V��$��o�9������\�9�O�_�c8`ి�e/���TQb��ǭ��/Ué��9]�F̰��uT��5]�
����Y�;��%���(���E�*O՘�`��r���R3�9j�2�]K�,��W�^���gV�lc�b�!����B z��K[�a�/��!�\�'F�G{����r�dlgu���0c���~a�1���^�.�t� #�t����p�OHz�8� �m�Y���9�����q�E���Q�ƪw�O1|�]���W�,
�'Z��@��0@�^��"��W4�tx�Y��FY�.�_�U:{�˴��p��K�?R�a�[b�O��#���AS�m�5�_��U�Qߑ �+��Ėt�=�QSL�6
�4k&Ӟr�;Ʉr\~�M�
�-���GG�D���V(z��?Eۅ�58���.�\�-`�˸��I��(�[��'
4l����+����CT�*�e/Z���Χ�ӘZ�F���;�LR�L�Aw�{vo>�T�F�(��f���S��V��hǙ�k��	m��jiE+%�-�D�@W�� �?��R`��p �,���s��c��x�8L�^��P���j�sũ���0}k�xE{| ^�����?v6��BA+-�!㑑>*VB��6�K=���OL����e�Q>WQ��(	K�M�����QR�����k`"�	`l���?~��5ȗ@e���#! �x����т��u���%��?g%�{��"���:�&��+J�/��M�5�r=?�u�0=�)'��I��j(�#U�J�2�>�\��:�Zǻ�����?-WufjY���y�hG�Z4^��aÆ��|
��)r�$�G8@�ϸUd��xVW��_����ʊ��RPP���x�hx1��f�ĮC<n��#��a)�RS*3*��E�O�{��O��fbE���|	�HC�d����ݸK��*��r"H��G�k���W6q�(v1�I9�=�L�ӿ�5t��0��8Y�}�Ob��Wk櫛��a����CB���ra���L��;Qo(+݉ti:�JKvW�5�v;S3eg���QD&��Z_�V�ks]��x����1���A����A��2�t�ӳ[��5�M�Wm�5����ـ���+k��!h���L�<%q�h��wA� �gt	^�����D(xR�W�K��k�(��tp]h�F��� ���.���x�f7�A!���^�4�u?��eܽ��|�
G-�8�|t�r7��i��� ��SNYI3M��9φN�X�z�Ҙm�Xx�D�.1�L*�'�p+1m,'�*\ i�1Rǳ����'5e�0VQ8�TFЗȐd��t�p9��7��⚱��j��bd�p�b��>�=�~Wj�E�j`]4
��IEX�T6 ؁e$�2m#v�u�?|	%���68�����?�ݢ�;���<��8��/1����hO�5q��S4���v˵��{�d��*�w���A��^G��-R ��!�
|̽����	�q۠NI�ŷ7����,�j��psջFj�k�"����U��%�+��.$��@��Q�;`L���e����D܅b���q������:8H��_�=�V���~���x�uzx� +	!�8�*]�L�y���w��\ �S_�}/���O@k�u)�ɮf��"�xi����s�I���C�g��F�ۺu��a�|d�tE)���qf�`�}�l�_���wg�>cL��}S*���������0\���@Q���K�3�� |f�E�a8��xx�T\&	p��qj�l_G��m�^�M�/�l�Iҫ�$:r	O�
�ğ(?zL����7'��X@�ѯ�DE�{*0N1w��C�օS���}�C�51^�ï�l�;Z��
�pZ?M��A�L��ΰ8 %�D:%�9��������K��0a���؞����P�D�[
�!R���1�04s\�f1eL(�[yOʹF��/�
R�l�d�G�w��*�'*w��b���	����W{�|E�8�L {�m�� �?�6�q���|�y��;�m��Q�C��
�|��=��)	�/������ �68tҘ%�֟��h�U�!k��2C5[g.U{x���s�_�焝��Q_���z��X��N����[���������{��L1͢��q{�|e�;��1�"r��U����[�O��'i+��qW��ַlz=_�N$&�d��� �n��e��~���_4��	�6��m����=s�N�����9�j���6j���S�[&�'�
L�zw�(�8nT�$4CU�j>#�΄�tF�m
�\a�d^Ťp(�Y�CW��Kʷ��5�,,vrWw-��(���z�I^$i��E.�������mH�2c&��Q�kJ�a���������^9�(Ǹ`O �A�!;ښfd^��q��K�R,!�{�� �$ݗ�:�0�ׁy�#z��C,L+��|ᵞmP��G�5�&�JU6^�����F��2�!����.�w��{VG���,��H�' UHR�*��r�).e�f+5Ois��\u�;2hf[*�=��@����v����Nr0}���-�!h;���?���ʿF/c�Uy1e!���v����8�[\p~����e�OnBpc�kA"�݈t��sN��fe<���-�V\杨)4�)���*D!�����'T��ĩm�bġ.)p��j�'���1�
9ƀ����[���#Y�⠣xѽ����"��ok�e�r��\>NӖR�!� @��ƷTm�nsI
�q�H��	 �ԡ0Y�91��).��r�ft|�Z����Y_���maz��(2�*߫M^-���&P��ƘyDM���`�����T�
�t����{�k�I�h�E�Hz�y�D�:�Y�ŕ00�Ο�T)k�w�RD#7��u��	 '���T A���-�.\y7�����_�B�����34"�*)�J�,�Q���Ŕ#�ݦ��%NBX��t��L0,� Nr��|4�J�E4�7���)k�ns����iCǿ���i�l�V���#�j�3୶h�4S̍����MǮ�4�i���; vf|���ǘ2f�m=9˵��u(e_��}��N���'�8J���i,#����U�w@�v��`�X����/Hw��1m�^�W�����=�JԀ�7�����±�Y �F<!\��^�3���Nì��Q�����Νg��*�tЅ|�/�0Q��x��]`�ܤ�,S
_O0}	1������Bg�`[���DQ͜?%�wP/����UZX�*�[J�wM/9��W�iei{~j�2��qw�E�C���}��X-���!��_��#w��ZE9���Iz/ھ�Ty���PGF
��]N�˝9��G�Z��cn�3�c*K&k�a9'.B�w�D��!K�w� t%�9I
�Y�������7��'�\Zô���Z�Y�Nlm��Z�E�#f{��2�Ae�Q)�v9��>��5��s����f|U�*�5��:t��WS ����-8� ��R�l���ը� o�/_ZÐ.�(�-�ÝG�Ť[����I��D�Q�.���r9)\�݅lYD��?2
2�EB)���r��?��u.���6��;�.A�����+3
T���.��6��t7��T��Mv"�QW��5V.�d|ê�������]��t�3�	7�jS����IT�	��5��>���DY$��-΢P{�by�h�|�)�/^<��ex���cѱiJ�-tVUE�|���P�8k|��Wa�^������>y��4�lK�׈���W�!��f&U5e6��B|�S���6������o�LZR)�N<�9o���ۂA��i8�P`�v���1θ�@䧭�O� �PQQ,}�_�/��B$����O�5����&�8������|^3Ѵ���d�=��h8��Q�ՉW�A��?�ｅ��:�ap��`�GNQ�)DyL<,�]3���"ڏ��_�y!̃(s�Z�x��2#�l������W<��J�
�}��6�u�3/=�#4��Įb@0����N)�^DSI/�Z��㑞1FQ��M'n������D����8�W�3��x�馶xQc<�PS\���
/kl�,�Hu�TGI��-C��+i�k�þlI-�r
p�cs<�H{Qt�6>������WA��t�R��>	
ﵾ4�
Գ��7���&��l+��a���|�S��/�t���{��v5��z:?��{���	\��^oi1�ʳ΄PZ��KQI�����`V�-+>���;��0]���pg�I��_�9���''*�q�?�Ӑ��B避��iUD������k�#3®+}{�CRI$Y�od%a'o����T=�q�;�>'ٗ�����h��{���^�'�)���a��8��BƮ$*tL�02�QI��R�j��m���]���:8�y� �qx���J�/'��#HE�g��&-�Yi����'�S*��+���ȢJj�k1G�&�"r���A�ca����O0���_���}&0�V�� eȗ��ʛk�A�|ެ�q|"�x<�x�wZ Fk\�Iy�tXL,��kh���eUD~��MT�AC��7�����:Q�P';����9��c7���ᶝ8�S�hE�[�!�sAW�K͵��a�W��������c�dE�@�,95)<`y+���<�B%�84�.<j�?@�z!��yo�������n��9���/�P�#b�������vĺ}��X��@�;K�W��q������g���(1�𳦶�1#���B2a���u��ԗI�3d��n��J]�Cݤ�A=)lmU�p�.ه�R����ܕTڅ(42�´��;#'j:���Di���5��y�ʧ}����Z��,i E���y��r���3>�R����: ��
��T����(N�٤���S<��CS����*�m����ի�����A��)�{\�7�ØJ�'O�G�k�f-�'�������J���Z1ȥ$���n�l)����F��7�9��|�qWQ¢z��8�����|��� iO�ho�IՑ��,ȯ������l����z�-�]غѮ鼫ֲ̠t9�Bw��]j.kT�h��T�%.���Wf��H�%�Os��(���?S���\7���]&"T�����#M�V���>�Y��͸�R?�/?�1�_���h����훐\k�e�*�!#��c�8��iee�2�TkZ*�D�&^k;�^�͋:VƩ`U���o���8�{5r��綒�'���%#���́!.3Ȍ;B�*̿��;����k��m���
���2q5��� �1�����D$�Ni���Iݎ~�MK`���؁�\:T���江5F���i���O�j8��z��$�:���ك5�n�����4�׆a�L�t��u܀�����t~�F�)0��ܑ����t\86fƼ�3�U	5a�M^|�#7���vB}�1�l�~p��ϚW|>���#i�o�#�gX�����&پ�%�F�s@����%���Yb�D�Hh�ԤY�06��?Тl7C�f(������'�(�k��՝[��EyC��07ȿ��7��<�D�q;=��L{!!����;��?�k��3���H��t�.�/��Cќ����_�q�g��cn���"m�c�[q�Iҗ(�K5�fn1�2�$BЫ(]� �\y��Lr��[��o�7�a�:�*GȂ�Q�:x>�%a�ф�dM7J�dn�&�"���'�� �Kh9�L�初�	��[bԻ���
<��U��&o3\Y�����]�4`9:���7p�BB��Oyҏj����Fhb�=>��(�x�˦�3��
�s�����2#�Mb�e��AD�'
�'-ޅJ����1�#������ �N?��PN��2��h��˷�6YmTD��Y��N�ɂ����	��v���@�;~v+�H�ĄZ]��c����/�U�'�ſ�q������d�$^�K�3�Tk�6.$�@�'��o�V���S��wx<�^�kŖ��T9��J˘hKc�a����͗�~b?V����ޢ��1&�����Yf�Jw����:,h�i���FH���<�ޏ�gu�O��?ѿ{��?�����9aՉ��!��j;�-����]X9�d*�b2b���|�C�t��MkB��F�!�k8Xkp���pc�4�F���gx�d�:���T�U�/A�g���F6{o&��"W;X�A ��<�N��͸-��A��Ŏ�5����>�bJϲ��&"y�}Ł���Ҷ�	i�5�����L��LEmy�~�O��,a�6�~�B�C5�>O5Yt�z�8�_�Un�zjESj"���}�e�J��?��C�e�D�r��O���tFV�k�e2,����yL���B=~)^0L�����E։g�6����f �0wA(A��0�B������Tg��k�6>-�N�u�Ӆ:���S�p��B�/ �6~tqp�<����D�#T���tl����mq���#�,�P��x�Ƃt��6+��8��%����w�+4��fHٮ9��B@L��و!�x@�2��#>�n�#���
sd/=_�-S-��R�4C��TF��ߡ�⨟Ǭt�����L܂N�J-�X�U�K�R���ˁbY�˛�UP�v�=��ݴT�Z�`:�w�%[�;�������`ߌs"T<&���K���ت��m}��<��ך�;���Nڃ��I�n���F�0l��*|~O����
o/���Gr(�Sf��!r=Ӕ��Ǧ�MI,�s���"�=��Μ��1����G��KIM~����.}g�%���û�dM]wyaH5d�D'4�t�[0�d�}̹G��0�7�9d,��s�Z�B�p�#(;₭��K<��%4��;��[�.݆���:��{L Y��ݛ`Đ�x��^;�U\��$��G:k�MP���c����ЉºV6)�D�C� �]36��Ԛ܏҇^� ���Q��mZ��g��bN��:��ӣ���M?�a�����t���6�� ���i맂U>ޜ���Z�����[�6�Z��پ�H�����P��вb���\GI��[�12'׉�U��"���p���)Νm�@B�$�&��y@�4��/t��M�t�F��3���ݿK2:�g�(NT��B�>��[����FZ���L� C���D�����pE��FS�N�QLΡ#Mp̤AG��u���.u)�^ɉ������.��ܒ^�w)�KH��e�g���e\`[��Xf���q�������Q�6ߜȜ*�	*��ӣ�w�N!�c�8/�U}�erƸ	8���Q�����/�F�W)��{�5Ajjr��uIN�Ylf��Ʌ'�<L_�����I�
������P���5��(�̾J
`�[�աd�]ҦW�9"EXP��)��qU��u=��B������n���K9n2�LO�i/���Jۊ�4��3Da�|�?N)�^R�L��yq�{M���D�v�Ы\R"��8�0�8P�w}H�o���4<f����B��*�0�r6�ƌ����G>���^k�YP[� '��*P�[���#n��	���^1���N�X�A���|qYء%���(����+�Vؘ��V�M�F� �<A5VS�����&����N�[����`��ɀ�v���u�Θp�7��0���Q�uKuK������D&��?<]EGșaq�O�CП�Z��v�n��_��C>�!�fǎ��d������z��Y�B���B��[�1ݶ+����0A�K! �4��S���2�U���Q�o��p�v&�=��_3?��q���RjH�G;*h���F�>2f?��bX�Kn�9�E���zmȦbAq�ᗳ[Ѥ*3X�>�+3#����!�$�J�l�O0x�X�.�m݇��@��w=AG\�&^�@ ���Th3<���b����+/�T�U�Yq+��z~eX+m' H$|�q�D!Џ�Փ�(��Q� ����,�ֶMݰ�n&᫃��mX=�kS�i�S���6���@���$C^+�TN�_�\0u�W��%h'�밽+V���\�̠y�˖�C�w����bk�^ʂ���9��<�O����1V��qD֞�9b��6��'�ǁ�n�d�k�鑇��	�hLo)�a`��nLv_��
�E*��^cQ�(j7�z
C�/Ŕ3�&X��'�T���%lo���a�!M��4Ȥ>+b�	�z⦆فvR�Q���]�:V����}��iN���{��J%���+[N�7�I�5�N�H��\�	D��� �i��!�s�j���w�A��F�����d��pc�2p���s�����-��x�g�YLЪ26�g���¶�j�s��,�ff:{��о��/>�S'���	��Q����>�Z""ШB��'�dq����+�%�h�+'���6��S��s�����Eh���=��۔£�^�ę?
��GX��u,W�r�����/H�w^ 3�w���c���z��~sg)q�ɏ1U��l�]���6Q

�#g-ZA���E�\����p��9����Q���o�_Nyk�MM��c�=�r��@�%%�B�6���<Kw�GWU���Wdu��d*�GO�iİ҇}���0�m,l���=5 l}"1X��AR��[�׹�����P����v�-�7�o��U�y���H�!��Zq	5��ډ���I�B�6�w\�vK��".���B��P��+��8�Y��2"BCt�'��SyEA�t��1��m������)�GX��n��������]����d���6���x�ܺ]�ЍY	���d�>W���qn���dE�j�h3\b}�[�,�i҅��h��ٽ$h[UO(0������\8������x�E�-}ǌ���ᚍYA��D7tUc���S �[ZO9Tt^��X;�e�x�Zމ.�d4����T`ǖ�	�r"P*P�Ea��V�>d�ҙ��~W����w�m r�'�C�B�YX��ě�v��v�J��O3����MHe
���|�q��痷`b�6�ԁ�(���p��%�'f��z��Z�54��M�OJǔ8f��l<9�_\BK���q�0��8r�2s �̅�dp_���}�aM%+%�i�v��������hG6�j���6+�d^��2|<����%B�.�����o����h���0�j�2cʵO-����k	����oz@�f=�]�׊��P�����fi��$��jK-KDd?�ULQU�6UMN�r�*�L�Ņ*�؏��rQ���5��t��QiVH��ٹ��hi��5�����%*Њ�������ҟ̌_U��s�8Vʔ:1�����
��:�;P��-�g&�3t򄻜h/���D� *7�I*nu��v�W_X�Q9T��%Y��8��0_�;��E�Avi�g���ҶRQ�@�U��s��R�?}�t'��t�:�9��$�LY0��YfުA���y3\��>��=����D��8Pzv����J<WG{/'Ô/Z�h����Jڤ���K2N��]��g�m����2��N .�����+m��˷�6<�����4k<!�V;T�X37�����e��61���˧)�<��HN�|y������!���Mp�rRM]N�I�r��/w�lQ+�dޭ鬸:��
���'=�t�M��8�����Qo�o�,�/a���;��F6)�(�s�#��%&#;�3S*��cZ����j�Q��"J\AʺӰ�S��g�3�>	��@~�I�� ȉ.@O�F$m=�#[�ƗƊ�	�خ�T���Ro=���Ή���y@-�Oީ4N������ Vhݷ�FR��w8���f��4����g�Qq@�]S�̱�@|0�U�o���������#Gx�6oq��S�7v�r�m����&����}��mĵURxn�`�eC%�pۆp�x���n%g:�"�y`l�Ҡc�ܗ���u�� �yWz��7�I2���x[�!{��`t��MXUajC�r�d�xt �{�Eu�Mk���R�?�[�	j�?�~�/��A\n�g�{���{Zv�K�=o���ܟ��_�6t�U�q-��������.���.�& :�����<����'�$d�Yr���-L�W�ژ�E�YU��'-���F)�&f�+c���Q?���Q8IS�Ⱦ�>��QF�`
azvH�z�C�,L�ͬ�)�6�,�[=^�����}���1�D�P�$. h)X�2������d0Ų:�x�͗� 0�Wr.�H�H
�y[6A �0�'��{�)�!�+�����8:��H��?��͘��5T���d�V��^<z�U�|�A���#-����շ~e�wui%�q�֏�1~ ��z\�.{�[&j�k5���F��6F�}q����UQx:����~ؖ�r��]�n�;&�JB�p���d��T�[�Ϣ@bT�(�A�G�8��s�ОC"ɂ�pw���_�y�-ܨ��O`ڏw?��,��ܲ�aLF|7�����5�����@EnBu����b�9_�Fh�(5�»���2���w�̺�ۊ镋�e��Y�A>c@}������4�y�Q��ݰ�hTݸ���=�����)˒���b��,�J|�|����G$�E=ݸ�	�hg�;����A/}��=).�y���6���6U���N�j.� ��;"�7��m��r]�*b�ဂ��6��(_$_[��(���~���jJ'��'��3�m|v4?�è`GI v�NW{�|p��{r�G�r
��u@�6&������&��4��#�3�B�:��0v1��5�C3\|s���zN�+�r��zN�ύ��h@5a����wv1dMI_�=ĺN��k������D��~����Sl�6Ԑ��@����᧪�g����!�ܨ���S�W�rތ�[l(���NҩWt��̵5�ȀS8l�̃���'�o�#j�����ޔw��"�Sx2���J�1�{Y�Tδ�s�K1z�8H��l>e���%w��/�ߙ7�����*?��g��ei�l��MI�O֒�h�n�m@�i6gJv�c�h��hh����5+F,�2���ys&.����[�Y�]�(�+K�A5OB����y%��Ƞ��;�wl��ɔ-��]���@A z�xez����;�=B�p8�uQ�k���
�!+Z�q�	JHe6}��P�b��8`�'�����>���`����.��v�ù����Й�s��p��ә�	F�0Z�� �*I�&x��''9哔_��yG��]3�T&x��\�ZfE2���Aq�v����u�&�簤Hޫ�{�w�~ϑ�R=X���懽o��>��m��/���[Z��%��T3z�`b�o)�:�3���1�H�C����R��&�������do�Y��]-y�}=(�YE@�0:��z����A�b���e6P���ݡ(�->?&�KIM�M0�D�wjfe���t���>���Kߌ�e�m�.��Cs�9�M��!E"���J�v�j�t�Bi��U&�S{&�����Q!�p��3�J����B���:����?|��MCg���
�X�]���C0W]�)��à*�&A��(���!8d~��h��R���(
��N#��ua��>��.�8�VƀiG5m��>u��7�*+�K�mbCC��2BrZr��[@�a�q���K�tV�&�8�p�*vDSE�c��b蘚那�͛	qOD�*���S�����\ҹ�o�;Ռw*"�\�,5�ve����$�0C�>�<d�U��,�֏�{3��3��1rUK��������{�F���j2���q
�=\c�������=˭�֔��;�;Ė4Չ��p&E�`ï���*<��22q��=�?r���v#�m�Z@WK�Y� ������t���C��In����ٍq�O�"�q;Ӡ}r����h;^�im,+�a�W�K��Ɛ��C��V/���p)3��I&";]�����ƻ�2��d��?
+y*��	;�r!
pbg,v��Qt��"O�5��}dtPm�I=��A�X���n~���o,i<�Q �?��ٛ�	�8�UQu�YQ��zbr��A*����P��8K���!����b�r;��ZO���C��.k� "����&�AH-�:-�k]Tإ`*�M��x�����f��M!#����zp�G����/Y�����8��>�f�jҳR����X�3�+99��Wϒ,k���o>Lj�iT���Qr���m
�L��/3M�S���"�����ܠG�539H���;��^9�R�����j�S�f)oy��/���Y�x�Ym����$'�L��	�>�s��$�s�&�W�A���Û��{Q6C&ԍ�;G�V��;�I�Zo���x��|3%]��c�?��oq�Tn�7�AK_�͔�� a&���A�$^ԗ��C�x�¯���rǯ�g\:p�����M�k7���Vڦ� '͆�:�H�O��R�]g��%�tM�����.w��)���(9�W�g}MW:�p�5�C�NB����p�������йE�����h�e�1�M����,tO�%�_����ڇ���X�s�E�HZ�t����{LU�#6qO�G��M���2��:,��	�+�u�g�bn\b��������S���j9������T��p��eQ��s�M��z�u�4��+��E���c��3�tC��ҭ��?���W,֔���-���~Llt;A0�xj��6��U"���B+ݔ�Hm�	,�`�W%�yOU�p��S�@�̂V?�6D7���۷ ���-��2���3�C�et�y��CAzI}��!�Sv��6];���K������R�޷_�>�^�,D�娂w�,���q���+�mgK��`�H����jh(��L�"~k��˃:Y�%�a\��¡�	�ʷ��C�è3JAQ��Q@�������)U��0o4 ��v���)�O�#LGƖ ���C�K�E�5�%�/���>,g� 	7|�/��T�c	V(�b�!A���䕴o��	�%q��\�D�5W���Q��<A�+����j����� ��UF��r�̭煉���Fs��Z��ѡ��b��SXT9�1
�Dt�3�h��,��E̼�b��'��	�ZR�U��Y�,/XLǈU�����#H�&L���x[�Pc��nN���q��HMu�*��yd:��D�Ri2�X��3��H��p��c.�(DK+�zۊ46+����x�`�rw�T蹝��>���e�a8���{� G��\Mn��J�֒��I����D�����w�t��3��~9_�)����Գ4.�fQ-�e�ǜ�u>�j^�3�@G�J,䋸YB�d�򯙱�]،
E�-rW��J>7��OU����h����|���
��V"�/�N��jp~��z����U�崌��⷗>�ʬ�Lp�%v.�/��蔷.�]��R2rG�i�a�1-�n;)[ZI�H�֡eRt<��236�a{��J8�<(jN5c� n_���w?�z���a��ᆚ(�����E	G ���|��{Ma�u�R����&�'45�,6�U��4��&���~��M�^��/n�
�w��7(e����XC�Zئ nh(��b�d{"��,	֨�ͅ�ϻΞ���t���I0���k̹�=������/˜'ֵ�\f�k���HWl/�	���u�XM��	v�@EM�58#[~o�d""����v,�Ȧ��������*�"ȳ�R +�zY7��X�>�G��	�z}����8�аHי	����m9��gO�ds�Z�@�xP�i�43����*���V��x����l#Ⱥ�5������0��{�\.$��c��}�.ή"�,��1w:;�����L����!��F�'��ww3��[���<a�S�1q%�T*Z�ߪ�1�U��Zz�g!ip8��l[����LW���#[�!�\�ޫqǩglþ��hn9�C�1��?味}m>�_��?P�?�!��b����0_QDb �
QJ&��*�N�K�Z[#��X����~��2���N�����T�kQE*���I1���� 2Yj�rK +�L�Ox�����
2�ŸU�Q����	�50{����Nj,�#ݡ�P�ŏ$���ݤ�9-�yz��>c�v�
��~���O�G�}C��-'�х ���ɖo��+�)��$���'ͅ{�V}�ц9��~b	N����J�r��QC�|e�L�6n�h��4�h@H���S��MRbQ���6�'�D+�J�>�:.���{6�nO�Cg{�$��0퐐��`l�E��Pr�ң
�5�H8Y�)��ת>א�'X�I�&�ڬ�����KF���!���MPsԐ/�� �ކG%�a.7��@[�w�$��U�Q�SA�p�?�>�8��`�D�Mz�e>�h->5�� �S*����?����:Y7|�����:f؟���#o�v2?���R 11�_`h��\y�@��5`�/��-'i ��g>�8�eop�Jk�����}W/]<P��g�6�N�Fp�s�T��s̬&Rl�F,]]�FZ�˵LÏI�$c����;]^����:��l�i����ݵ�2���z�3'��VĢӑ��S��yy��k��Jf�׽XB����]�.�p:ŗ��t��20F㺽rr���7���x� ��;{i��dC�����(Yc��������
����82�z���»B���v\�$+W�iX����V:r��T�>n�[��̘ؔ�2v�Ι������!U=�7�rMZ�w��MG`��1e7����2�b	�����5�b,���_'��_T�/U��ǊO,�v�.���(���Йx���� ~�q�m����e�Г=��m_����D�(��&��m1M�	yB �m����<䘦�c�SG{,�CJ�/۫w`��.�F�^{��`O������:�"�(�蠑h�A��F�l���y��p�u�K�֨��L��R3<�|�am����H\�T�[�f�ot�wFUJْ��f�
}<�Il���Q��!_W��G�`��9��%r~��4�΁�סN·��6���4����?bo�������z�/6�oR�e��B����3����ԣg/`6��b�5�s3�V���c�(k���D�t������3��9��Ư2���d���"��]�ԁEr4��5U�q�����p/�A�V����ۍ�)(<� N@��Ԫ#�u���΅�i5�ʾ�2�<������NG�QȈ�iM��X��y`��fF&�E}K�a+?vc�'��3��D^�AA������z�ΙIY�794?�I��y�-i�9�<xP�j����� �؈�@��R��"�H��3��t$�g{s�2og�E%�!9�e�`��{���T�@��3�M���k%�3Uʱ�3SQ~Γ3�?zS����<F��(m�ǌ��iT�fl���u�/��S�+\}AF�N�°]�C����9nA�2��h7���z]r�O��"�1Z**m]��gN���@ᲗS�}����� ����%�=������b&d3b��u�� S�ei:a�ز���+��OȎ�㖸K�����_�1���g?�n�*l��,Q0���8�|��Rd�$h\�d��-�m������2̈́��p��
�O�Z�&Q�I��7689�ɢ:*��8����i@�J;��cv*q�-�А����u�jڢV�B�VP�,�dX�Xy̞!�����cA���,5��C�����>�Y�$�^���g����,��D�Y�+��0�'/˶N��}P{���I�n��)�	���Lv�-��čN,�=tH �4;�u��������m��<�٬��7;h��w�Al5hM�q\H�6y}��Z�ݱ��p�8K��Ȧ��)Cl�����%1����ϒ�Lwj���I_m��KJ�;#��=�O��Æ�:<6%%[?�3����6.s[���Md��p^1^�8��-���'2��/�dًN*8���Yh�Zr���3�H��]�:�ȫ��F�AWK�C��B��=��WW��8a T��FsGj�c���mQ7�������9Rt��%�Ǭ8�K/����<h�&�'**�^Ҥ"m�_L��3� ��K*:Q����۶��~�Ź����D6Uj�;�L�NR��w���*���k�c�&n����"�}�ŕ�)��a��GW��Ɯ�k,�[���+SiԍjC! `�<��D�X;N��"ɲ�k�O ���W��+��)]���)�Ua���&l`�ɂ(]�P���=c�r��
n�ر.&�@�aL����ĸI��biWk��SϘI�<(�W�z��:.�&��u��JEe{pa��/��tL�D�GN�����#ש���#D�q�����w��N����T���A��R��������fQ����{��L��Դ+3f雸Qj��I��\}��X�G-����3�Ԙ�x,���V,�Bh��`���S,wK�C���R}=����H5�\�?J�	zY˝gZ�Q纝�7����1ItQ繹k呸�1�����;���v��&s��L8���ܔ�]ltC��r���	�_s���jLI�ē�T-��(z�d���jޏ������p��>o�Z�މ�:˔�l5,{"zT%Ì�3qP	㪹sV�c	0��@��lt¦�&8�:��T��U���_�bp����N�n���EVA�3� ���L��<�}�#-�:I5�>Ж{�� ����õsFR�}.�n?ԖQ5�S՛�^�K��:�	Z�X"��79���sƌ���R�����"{v?z?h\Lzq�M�����Q2��̏�i���ek9w���T�!���4���_փcY��\�,ݻ��ߴ]��~��=�!Нũ�9$$q����R�f�RI��C3M�o<�`j�yB<���l�'炟��$�)���w�ـ= �������m���l$��1�@Ѩ�W�֨��n]p�=��ܬE� �LV���_��?��鳡��Sm!k�����_ZПI�(	�)��~�V3��e8�ᯕ�>k�Q����N>	��n�I�aM���]���N"����хw�|�D�Wz�+RH#1#Bmx<��l,�"����w]��)J�?ꩭӦ���>
����B|�B�dY��$�����E&���b̖֗
���1�&+`ݬ�M}�O���la�E�rEC/�<� 7+#4V�N����C�O;j�z����_�ƭVn�T)c�~��*Z��1foXHg����"�.�pT�S�s�@��ڽ�9��C��`?CcP��m��G��ց�ɤmOs�F�.J5�j]�^���}��6d(�$�N=S	IS������]��߾;*`�Vӂv@D��Y���!��@�����;���5&=&*'p1���p�.u>I���_Iv�8JTL��z���Y�*]�K]������}�*r�l,��/�7��N�L�m,؍O�[�S��78���������/��L���x[�V|�6s���>�S��:CM}�~�[���so@U=�κ�<���x�I���>]bh1Ŀl��ĥ�\�w-�;�r�-g�|̆�����]�9z�GB|}zC�J�tI'cS�����	�"{E�����4z��:R�w�{u�H���̠δ�a��^�14�اϬ�nH;��U�X�C����+�1�z}����S�-�~M?���BZ���i˓�n�F��W"�����7|�s?]��K"%w�6�$��AW�QPe�?�1�xl�mr餜�̇�WJ� >b�w�K��<x����$N��Ǿ�a������7YYX%��훁��$|��5궛���h�IHx1�tD h�">��RX���3��4��j6��<`�*�/K��EB�����V��Sv[�����]��AV��K&�r�M�,�U¦?�[����*3>ScH�)~�����I�BJy$�D����jEݏ7�_��!}�L�*�Q�$���yK ���N�N�2��6W�X�|��Qzc��/a���2<�_d� F�UːkI���X���B2��Gg�cfȚ�"�����>����J,����y��0kX��bׯz�j�3s�@�n�a�ޘ!D�Y%_f���]�!��c�O�M���$��_I�X;K��]��-�Wa�x��wg�o~�.
AU{��/���u#³ ~v��0Ĝw�����C�I�����&g���Mj���nf8v�/�Zd6�4��V���OB�z������#XP��;n�a+�lG���������k�/+�zv_��J$�A3l�\/L�Fq$,��I�)p7�)�Ox���X�dR*�B[�|q��P�}�_-��a&�'�{�nB돰��5l��DDD�`��,m��z���>.��v4��+̲f��4��	=I�Q���v���,��x� ���z4z�o�~�̓ 6��v�6��#}��X����{�k\f�v�s�6<O�5��ʷ�s� !J�7i����
J_�w
q.�bo�3�����X����-�_n��3�}@�l��}�m�v_v��e������8�(R	��`r}G�v���x��b;-U*BE�d�����>ϖ�g2ک�ݥX=z��~���0LnkG�����{}u�i1<��cKDD-Zp�L�\6`�`��uyn��3ߐՄ\��mxj��A���>~|��@��/�z�X��^�b�ͭ{,�^���V�Hʵz2��j��V����������B8>��"Ut,Q9��i}ܩ�8_6eז$�4��?m}��,�]Th؜�}x��\�1�����C�_C��2�_��ʶ�x�n��m�I�pJs@�+Ǿ2�4�$������"r�j5�d�X��B]Z.5٫+�R��B�;�A^���ިM��DŴ��qjU`�����O������,�5н�ݟ�0&��؇��#��lk����=!��Tc'b�ۋB-VGʜ����,hSɉ�}���`ƨC)���Mw���^���o��e�]�==��+ܚ�E����1
���u�A]F�վ��S|�6���.m�+7g/iU#��?x>O�\�x�|��6g"F��P
���Х�4�*�����.1���\I��լ7���Ao�W'=�J/.�2~ѮQ|#)���!����J��s;Qo�/��|�˙Z�o�$��6+��·�g?�:FʔaL�K$�?p��8X���[�<�n�0�Ox�d���+5��s�_���@h(�J��d���W�u�����*��tfЀ5�>58� �ZΛ�ڳ˔�D�N@#�Ķ�!B(����ֳ�5�4PY�K-���bm���J�C,��8�����Ӏ����Lyw8�f_�Ä�*]���Ï*�#��_'D=���5�jU��T5MK=��2�kt��=N�Z>�TՌ�֠#>�_��"TA�x
S{�Kי���y�YծA,o]���yK�j�H������x\{�{��H�`�A�ϟ�<ˑ�8:M[��	�zؖѡ}M�!�2E0�a@�*s��P��7�1뢇
�Q��Ȓl��+
����߁���8��A���w�fH��c����!�ߐ��}P�^�`B�|�C�u� x�'�6��ܨy6Y8�,��*��S^vڀ5J���g2����g��]Ս�elV̫�'wj�47<��4i�6��^�X6z��-M��M�%S���ݳѡ���q���W�@n㖝���T��U��o/�,�]5�K������ĸB��P9<aUmވ�ȃ\{����柙�Fw$�{4:~����Y�:NN[�=�8^5ni�^$�y��rb�1:M�
h,+k�����.�?�!�G��7��跣.�4M�rчD�nm�XS{�0����!��MW���Y�^�^���c���z����x���9����-�m��i?ˮKH��կJ��`�,N�,�8��,#����Ӧ,I�f����ᰔ��a�:j�lM\*��+�8K�q��6M�,7���Pk�,���b��4�/g`�Ȁ��K��G��R�`<��wk���Y��8[h��2�Z������q��:�]-��E&G�ZR�nd���~�b�ӏ���XhЃ�'�b�@��ӎ������8t$�:��.8_�N�y�r0���7-��g=�����/>4tq�tY�3�'����g�B��[uu�E�ɣ�7��~�<���OO��$wU^���Q0ҳ�*J<�0�X�r�K�|#�Q��W-h�+DY��� 9i;�q�W_�S�ַ��.���/�F9 �Hj��6�Y[|�M��_]� 	�Bg��T�;b�ŘF h�Z�u�/ʆ5�#��gߢ@ۧ^�j_Y�w<%����ֱ�8DyE�"FFLYI������~�22�������R!�݂+�2e���	��T�5D������ֲ�x��Z���+$�q�#���bP�8D�G���_x�[�#�K���¯��{��l�y���F�#������ٖb/?�ܱ���4����xr5�Ђ"��
,��M$����<t8ͭA���AI��y���h)�H2tD��{*�����,W�S��MU}�+n��s�gV��#����ݶ�p��rCq�(��y��x
�2s�j�.�lu��@��nl���Un6�:Kz�np����7��tk)T� <l|j[=���`,��IO��i��δS�2Y�� fY|n�)�6漐�m�~i���^�4_�5{;>G3#TR�}嚑�KɯT��1��s�l��#���t.FE�WW�Wc��]l`T�е����b�a+��.��1R���F=HQ[����Q`^^7�����pz���l���L)0l3j_X佥 5[�ޢ��q�(�6�b��Q\�xrQy���Υ6m�U�@٬��H�\zU?~j-X�Fa��˄���#��iy!ؔ�WL`���=�o1Q�k�Ϊ,��,���\����BGo���Ő����v?-P������*u�wĚ� q'z���,,����6R��C��z��6���CIt
m�W#e�����C^B���O
,g�<6��ԕ���Dlu��_�S+��y��X8 ��SA�P����l!fG�zznܽ�V*�o��^�9�K[�N��&�D(F�B9}�C�4����&�b�o����G������v�O�h{Ȅ��8���ˢ��O�ѡ�YԵ�	x��8��@��a
�_�K�*7����Sl	�%��tm�况�Q)a���T6���5�͖��,X�}
���-�gЏ.�5�A3/U:N�?��]Z���z�/I�^�nbj�;��&��k&M�z��4��Oti�H��Ќ�l[��)m:���̂xg��y\���jk(��6W� ���4N����A|+�*R'�٫��}m��>���e��`i�k���bd��U�����/���M�v�/��-pW~�k�h���k��I3[����7+q���j~�C��Q0+vz�9ȹF�gk1��".��7WS��n�䱭mhDĸ.�Y����.�
FL%��?�x�[�HG<�u5�$ے�P�]"̋�uT��F:=H�'˜�_�����eӄ��5R�\�L�IG���S�9Jya�uc�[EK�����7`��c��J��>�$��ޮ2��nG�Չ`DZ�+��F�ɮ.��FFWw�\��%�*�9#I�H�@���2��ȓ���y� 2R�-�K���G�W��a�~�K3	�%`�(u���g^t��8���3ϒ�WP�C�
.���:�U��}����S'i��H�}�IH_�ptد��������X�2��W���w �4Z#����ֶ�40��8��v;e�	dG?�|~C�/���l�P@{�����P�,�L���Į��I
��"�>�Pύ�B���}���͛Y�d7gu:1L�<kE�9"���}ڽc�r0������d��h�>*xT�+�#�)�Z@���%,F��0i©]7Vd8��hѱ�o>b6&�h�J��w0v�����1����� ���@xk_d��8�@6�/cG:B��|xI
��|]ڳ*�A�A�����W�d���x�83�	 /���ٽ��ǥ��ů@h�MD �e�v�l��N��rWx�b�	���,�-�����)�򞥌2m��a�H�=�!����_U"T�T��_�6+3w��������9h�!�j�����;Q>W���n��yIN�a�jQz��^������T!��.qJ��7��#�/�M�E���$/�F�{�ߠ��f5�c� k�Aо1v\��Sk��D߁R�}�Y�� ���Igq?��&�J��ⷻ��cE3)3 M�;��u+4�Ho� �&��|:�]�v��ض��	%ȩ�2��^y�t�]~ȫ�9|Pټ0�5^�����?�,�VRn%���V�,�33r\�.���̔���^�#�<����d_8N�E�P�G�x,��L��D�xK
�9����QRn�&�||!B۝O�y�d�"���l�rA��>�b�Gׂ
"��n�����W�T?�T�ܧ���.B#�^t�\����6�)@��wrL�F�G��0y5]��t}6�W7W�͸(��u�@Ƣ���]�_!��r2%�G)c��L��x�*T�S�`��	¾���ib���д��M��+�����,�	����Ο��ثƶ/0h�uEeݧYR	g�i����	:��,QW��k������!������~��yv��o~��o�
��qB�!�,y��ݸ�{����\�;S`0�,va/��ej.���v�������ō��: �y�̏�z�SFT�D�켆{R�)�����b��̴�{�r!}~�]}�PLf�ND���9�q�,+���:эd_�������Y|�����H�k\�l�*�2� ��8f�8�Hzp~��=���7�|L��2)I������z��y��6�@�vL�9���j6����s�-Se��&Sv�����TLdj'�. w��D��2����+�#����W�Za^�C��� ��K3����Hz��:ņ������(�o2�<l���WF�#����3�B��V�bZ,B�-�|�9~5���笁���ǌ�3�29��LNM93�h��\>�X~OrhO�eoV������sg���4���jU��OD�J�bw�)Uf��#W��M�	��Eܼ�T|�Y��a �J&�r�c��ʀM�&�h���NKo%A%ȇ9������S�yz3b��YMدiN�;��A��C�;��d���r(�2GA�%�␿�b>�lfsu3����c��#�� 3ͯ�����lY}>�Ϫ"������
k���WV���r���K8�])3	D��B=�0�cz�Ua�/���ʄ8V��p�D���A�=E
X�+oa=�e��f�5nq�"�3�e�8�oA�"S������#�^�?����7���k��D�)�n��=e���b�=U2ݣ���RB�+n'�v�>1���i��T�0ZM�.{�ޜU�K�_Փ��B?;/�.�<�1wy���F�.B	�<
�G�<or�
f5��V�uFF���T�L����]���Z��fbB��o�̎v6=��$���ͷ��m�ĸ	���9��kI�<KЪ��2�VYV~�ߠ&i����i��2���I!�|>�ܕ�pO�T1M��h҅&XW��͢dF�@��^kY��#`e�#�����z��E5uN�u�PO]���(	�-�Ԃ.�=��5@�P�o��:���LT����H���"%D�+�%{��-^s�D��9�Љ7Q��jEg���^����ނ���Y�(���{��,�_噀6�����I��"!�V�q���zfw�u�%�ZSk�3��J�{���d�:����uTH��h��P���* �0�)�P�C�'z94�i]�����7���7��iJ���Q��I\����*m�zm"�
~"Q�崙ɝ����H����ær��Y�ĭV��>d"H�*��e��X�5> ��\��H�]SBE��&����g����i�d��,�6v������?�`��gs�5���!WS���>BА9�0�i�+���@���Yh� `0�Y�_H#W�2��I�IwYe�bI���iMX;�D ?xb��b(3���P=����۞3�x���Hb\�f:�V�@{�)S�XY�D#P�<Á��ϓ����~�ay�>�{7��%jc�L��q�G�,�α�e�S=d�AU�F�����Ԯk� ~�(l�Х��z���C�9��#��ș��,��
�t�y�I)��}j\���2e� 98i�Z̕�M)(mi�
~��ٸg�66��� WF^�4� ̀A�'��p2~����J��JB;j�*��9%[U�~u����7�/��W$2��^I�.�"������h��C޴���C�L���bEH���}[��d�xp��T���4#
A(G&U�6��7�,��j ���ʖ���Jz��8��&�w�xfT\t6Q�\{�i�6��<t$�bC�ݯ����$ڄp��F �E4..9������I��O+nb}A�c�::Ho�Rrĭb2`^�Ҁ�<�!�~�&�0I���_�?����ƞw۠�Pd�T D���+K��v�����b H�{ݸ�-U��I��t�3a��Փ��}MEC��@稺��$��^Ba�8 �d3�4Oy3�8�HV���#}K.�D}��^*��J����47�64���y�J*K�}�gDP��������N���m�|�Ȕ[q�&��˗�j�y�t{�Y��q�h����h��4�"_�M��[��'�!~@᤼����i�G��}�V�Z������ 0Uԇ������3��C'��[�U�t��ދ���n�2����_�w�1��[X������JnZ�e�sJ�=�#,��:�|��
��b����9	r�#��^O|ޮ+�뎜2(��UNw �j5�iݾv�w�#*I�M���;��>��g���n�C��pǋ���)�ԕ!:��*��H�Bq��?�ʣ��7��hy�N�~�]��!����<6�P�Jf�ne�كP��������ʹ��`#��䄧8��[�߹��$�0�7��S���gB�R�&�I���4�,b��=v�~e]bb���z�ȁٜ~�
��J�|��؃�[�1�S�=�Y�(~��W<Y��@pS�2ܜ�V�l
�?��2��x�M�NSi=кP���=M-L6��5��#c]�3Ҥ�����ڧ�Qя��E]������QK�,����5Tk$w4�Y.�С�3#
н�J�7S�d�:���VM)�[�Ϩᖒ��4����ش���8:�fQ�
+��x|��@]�u/�^���L'��Zr
 �������4Kn�~��ߕu^E��C�Ģ�P7��*��&Q�_��&�������6ɔ�Z}\	���R�^C��)A�V�E(���D�-H��Ϭ��7�`Xj7����+X��*3�t!�
X"���C��������ɧ��ԅ�Z)D��Z,bp�T����%_��d�����b+��gѱ��/�l;�!������3Mey,��v��T��T	�D� z+
�(�?9��
B*@���P�D���F,8�����df�a�K����94V'�0NEN�<@d��G(��1�oT]�^��ݐ�ؠ��6?N�<� x����L.>#i��^!/�B�,��
LC��&�|��W<W�t�H���K�!�i���RWa.��0���>��2L3K�Hx�f1��D�@��;��M$��ۈkڜ`i5�F��I8�?p_3�}^I6�nk�YWhFT����.������'W�-����['2omU�����W��z eTwv�uUtN��^�x�wP���lV�����35�gl��Y�a��y2��W�"��c�#�ܜ�$y;}����i�)Alݨ���^��5Β���i��G��5	!��Oc�2�nP��}�	�nPҏ��w�m^�UZ*�ϵ4mX�<�w�80����C�K�G1d�j��'Q_�>*jr^0��-���^��I��M����ӻ�sg�q��T �y=��n�"��]9�:�59S�ʒ�g������tFO���b���}f5g�euX��)��k� W���)+8�*��#M�-��k�����ȹ�{�KDp�~��k.��,׽�K��o�*��7�|��+�},�	!�4a>��4Z�I{�(�L;�Z�д~&K�1�b����y�L�
b��Pަ�R�H-��	������4%��R�\�YAז����u�+��D�3B]��J	� ����Jg+X���� 	VF���T��%A-��e�l�.���g��Q�M��`�>\�Yh���O���Z�_pye^i����;��*�ϡM��ޓ���Ӌ}�l7�r��F����xNz���|�r������ C�Q/0�0�t�2��O����?��J=d���6.�9�왎M�͡{n O-ۡ*�3>B������c�滷��Y{��w3L����d/@�m{�;p�����#b n���ka�����즂K��2OU���c8Tz�ք�76ߧ��rv�X(U�Z]���
�I��B����g���\L�U �Se����5}��⚻�����cTF��Y�;�'����+����������i�3�����[�y���4l�~�B�|Fּ�_M�����E52/-+ۤ�+���k���=y~g�!2U�L�l�IN��%&�[b�"�~y���~b ������nw�Bx�íkH�����s�@�.��K,��ɰ�E��+��
v}@�\�{�.I��/׮~�T4����v��9N�i?�B�9��"�t*���,[���h������OC���J�P�������D��8�kׅh����wܘ'�FDS�&�Y�2R)�!����w��1o}���8m�O6�D<��Ӷ���+��������	��Hw�8����69�?�!�-�lK/�vXRQ}��~�j�hL�_�[C-�%
�{P��@�l�3�B���v��|#�
Rn4��9 (�W�c�c	A���@�k�#����@��]��|�|�Q2�_o��*?��%����Iq�(�{4r%�ɰӦC]j�{r�-%Ԁ�]�}A�8����v;�l*���1�q���F�C�o����RY���#�>����}�������-��.��N�[ɕ��L�5���P
��UZ��=~ر�wWg��2�j�jc�R��x�ҞZ{ros̸ʔohX�{Ho�Q����W �����Fp��񀕨/�C�M����/�t���a��%;�x�Yk��H-�g֓R�O/G����Lj�����{��j�·2o�7l�c�J���L�$)p��z���|��2�7��24'
��F��ح�P�a/�/�h}S'�]����yi�ÏU��� @j�8!!�9R����^+���mXY� �:OL)�� ��DN@e��߂s�p?�G�w����Cs���;1�X���ۂ÷��u�R�3:�Я�����X�4=��?-oq���m�Eƛ�3@!LL�/;'U��,��2o�zp�}�6\u��F{��a�8{	ʄ�12��k[&@HJ���9���uBq]'Z5�<�BX�l�m~��ϛl�̹BE�is�sBM����g��G>pg����u�m�Y�2/";��M#p��72��A�h�n�nHIK�
��o�����rZ$�E���g�-�Y�H�p�Ai
% Jc=�G���������{͕(��Ǳ}i�L^~vR[&u"��$����x>V��w2y����߸,�}`��S�)t���F�4P�(�eW�?�Zw��n�1�)�Ȏd:e�&���lP{�e-$�� O����`�����7OC4-d`X�q��g﷑�����\��v ��]�!F����ie2���f�C��(=�_�l�8��[����.���8`=�!4r��d���-/崹�6�.p3��W	�Q����Y�������x��v��3�i�19V���f��� �>wfϟ��1�$ '�q+=5�E�]� �`�o巛F�kk��=��fG�0c�AA�����_��:(r4A��z����f������~�_�'��ܚ7s�X�|�y1j��������Z)9篘�e|ch�}�:0��Ye5�<�S�|���볺ǙNK�o����
v`{}RF���/bq�.1ǵ���:�?svF�I*��df/�s���o{0��!ݧp5��^`�|YZ���?����C�oD�,(���^qk�u�t���� Mf�Ӡ=�朱,~� ^�xeqB��u�eL�	�X�⒅˪�z��wJ�\���rI���!s|��X��cjH(���`3��~��C�!8%�����R�d�2NؔUYk��vHo�	�L	H��'B/��$.��[���cf���0y���؇�m"g�9j@�BCS����\j� ��8��$!3R�f؆�m�{e�)�x�l�.O|k-5v46���ӧ7\�)2dЀ5����ٮl�QǇA(s��nw��\Ɲ��s9'2��_�i�%4��4
�3d��>�d8P˶`k�/P<4$����X�1��eh��}���X�vÈ��*
L|�:n�$���<cÐ^B4�J������ia�]&�蚹{=��=*�>�r���4�5Eɩ��������C�%�@Ӝ^�w�p&v��H��2�V�@&cBaZ��V�	C]S��d�
��5K:
�1����G	G�*&}|�8��u����߶�YȔSk� i�M��I�����^O��3���ap��t ��S�8p���a��n
ej�:���p���>�]�D`�_�v�f��]�6��]p�bh��]���SF�[��/�H�m��;���=��j	&���iէfT�8���U�tf�4�\�U1��k;�]?̤��z~���߾Q���o�Z�`�u���JP��Pn�@�Gy/�q~�9�l H:�!���mf�	��R�n���JA� {�yE����u[Xu���#X+��/C�(�������-����G���U�6T���Ek��մ� �
���i�q$`YD�'+����̀������|\���y�H�V5�ux�mϼ<x��Z���:&�+��v�d��B	z.���\^',�S�)�JZ�p��=\_:�,�L�[��˚0��6����i�.k+v���o��.,Ae�XWjX?lq,]1>�תU��pm��2z�2{K���g�9
߶�E5_�[���[��q�^�+Y%��)�tW���?�k��N�4�j���sn����w8�)
t�fN���C��<��h��N	�J`�5R�ޘ\��d�݉9�~ �������V˚��3�G"���9����q��^�pw������'Б���BO���f��^Fδ��ݡ�$�Y�sou6� v�[���ܿ��}�_�����|:c�)�!��#x����nm}T�ƃ?㺎*=Ll�$հ�:�^��l���R��~a9u���w� v����O~�iɫ�7�J6|sz�3��B���A����H���j���+z�t�xY�����|�̤G<�`O����ʇ֔9���NFB!T�OO�����^��p��/U�9�n�<�gi��@S���]�,����Am�]�ZWH%`�W�i��a�ǆ��A�!�1N���mX󚣻�Q��<X-F�*�}u���x��F�X�w�>W���0�
��K�6%��pI��+���T��b ��BT��u.�����#��W����3�Cv�M~��*dlΡ��t����en����xtkKܞF4̛��V�*\RgCw�7`w!�遌��2���qX�<��PZ_+�d�sr �Vd��G��&
��_Z��R���ME�;*�?v�l Cf��yi���r�ߌ�~l`�H�m���ۆ4j��!x�_��&h�y�VQ�u�G7���gƾ��!v.|hR��o�X/�i��h��)N0Jl�ȼV���a�(�*I�1��T7�P�y?�8|c������_=��6�|/�v�D����$:,��p�X)u�uG�5}
ce�a5�������cF�Ǖ���i��p{_̽3�Q�P���jt|�R;����7Ss��ct���M��ߵ�G��h����;з	�g9�H�� c,{/��ّn#���W��'����G*���b��2���꺞IO0��2XC���c��q��IKO��%IB_��eĴ��ԁ��K�7�^�!��5f~z��N���;�v�=g�ԹM�k�Xz��u�I�>�����^�Ҏt���m@r�,�����Y� +�dq�_K?!g��i��J�;��8c(��bt���H<D���}�.QQ7Ϋ�����x��"G�)z���=;Q����
����m��ik�/��%/�P��C��!�
״���Z/��R�H�fE=kmO$W2.��k�y�8{�#��ˡ½4`��0Y����s�O��<�ȝU�e��M��C9U��fdv��1vU3�s���t��9G�kF��q��w�pL;c��n� [O�ޑƇOc�3�%zo��K�l��xQ?��;�n/J���!�+f/�bI�wx��y�0Z<�d�Q��I���BV��䊭 TІ=	�'����&��<L��R�qi'ɽqVk��Ö�sL���ǃ'�a����Ց&q�{3�S�.2K1r� ���¾Ú��y�����@Aؕ�D�VS� ���-���f}�����̝��1<3,�Bt��P2kٲN��N�(Q!�>K�J+�$����k��V190/��#pI�6��]�ȯ�����*F���'@r�U�����3�lڐ���7��]�!F�p������>��Gm�;CIkU�h\�;��@�=����J�L(�e��[�$��Z���Yc����������b�9<�bk@.�z	3��H}�񟫉ܥ�"��)��ΈY��j�7p����O�����:� �8|w��r��l��ԝ����8���"�pg��FF�TNn�vڙK؜c,)u�����e����>�o#m�}|K�qn���~7n�A�o��W�_��L� ��v��G0�QޞJS��-���[�����O2/׳�?�?.�S5[�_�����m��P��a> d�xϿ�8ky�3�����w�� :�/�p�w��{�ޣ����B�z�rd/N(?*�ż؈�<��Ѭ^)��@]�*͸�q8�Bi�v.c���У�T��Eߡђ��.N�+�F��ݥ4'C(j&�QNR?j��m�`���6�e�}>q�8S�N0���j��w^�%hi���G?���iLf���M��|�x�혡��޹�s)�H�K�Au/a���gvŰ��f,,�x�_?��w'kAT����h;����p�R��R�̂\�ŷϡ��S�wX��?�����ۮF����1��>a�l4I�Z���f~ pf>O�����F��x���F�&���<J�����ieГ�z�sY���Ģ� K�T 8��Xz�Y�����*(��}�߬WY���tO�Yf3ֳL�|жh����L:�)uW�\{�d���]�`�ͮ7cEXL�����Q���`-}� Fy�r�%nC���E��^��3�;�:���s�o-P0M�n�Ν<���#�Vz�<лB���0pY��i��D��{�݊���/jÉ��S���z����5޶���ٙ:Iz��ē�,+��� ����&��q0���_��X���Pz��ނ*�ā 0u8�ɉ�RW����^�ɢ�(�y�aNi�n��Dp�[t��B�t� �n2RѫI��[D4n$`��%��<7���+Cvn���5�!۩�(~��I[x�K$�Vc%��D~EoL�e���ǋ��*�,��\�[��7M���Y/��S'�ד�^�#|��"`ͮ#�>���6�DEP�z�cy: ��-i�}��<���q����b<+�g��%h���|��0Q�� �t֨��~:֍�s� �cߩL&�P�0єq��c�1��м`�������W>0��@ih6������f/����u���z�y���ˢW!g�Z�Lum*�E�(y�E�G0�Q�a(�h�CCs%�ٳ��Ӭ����Jt�����,�w?�t�d�S��Ϛ�+1�f���*m��y�4�hvER7f5�W�������rl ۊ=�.rl��ݬP[GE�佋&�[u���L5�ݫ"_c�l�'�I.�ݏ�A8�[���n�Q3o\.�W&����>f�-G����o���[�&a,�;�K{cE[�{e����s��Z, '��]8�_Xr���\��ɷ�8�1�|PF�cY_#@7��c��:��i�HH�סTA�a���f(���㍠K�O��[S������bG�T�"��ǎ�h�W�b�)F��gI��1��5�#�Ą�iN�y�E �V>���_*_�p�T��`��)����rǤ��Ŗ��� �d>0�.dd,�8:{p[H>G*���e�-֍V���U_����m��::8W�h�K��XFK��b���#�z�Df'Ì���V�.V"�)�b5i�}�l�.W��T�4����ݼ�f�u��.m���4��9�j�H}�ߛ%[v6����mA�M���S�G�8O�D��oX��g��"���:͏T&6_��c���8����/6�M6��m$�^I.J�S)�����6�e�S�<M/R�'&XjG�tﭶvv������녚}/����Ĥ4��99��)'2`�� 8{ކh�W�4Abȃ풟���T��n�0$��(nX��,"��Ř��������8а��L��UHέ�K�N���F�I�Wi�~4ٜ.eS��Z\�ˁ�|���h�^{w�wj��խ��h�iiPwԫi�Ch'h�� K�I{�|l0�NB�T�@��r�ˏ
��L*U��T/��o�Ħ�~���^�1۝��x�؍��k�)�6i���v5?���d0�[�CCi:(��;u��f2��]L�y� Zw�d�N��dw��Z������Z���[CR�����u�S���FF��=_�ܪf���>�� m�;}[�YQ~�(���r��G��)��z�Ոk�ǉMčKE;�[�t�L�'�E7oCVy=�U��Z��I��!�>��'p�c�s����
(�kaX��h�ΫkL֢|�W��W̩.�.��8?QD�v��
>�h�\&�ww+-�^�s%�O��I %֖!@RA��NT0�1��9�S����×�}��	e�M����Y%�U mh4�$��M�$�,�z+šh?�+T��5i��L9�q��~n'�cި�*�"ɖ>ؘ�(�������+x�2�#���hp8�M�	C�3h\x-�$�s�� �̇�	�s�z��)��z�w$���4%���҈�`c{u��C��d�D2�<�#�]�$����S`���_���s3>%3	~z��T���#������${e.R���J���8��\5��nׄ�~��W�_�-v�����]����Y��j���C��ܔ���K�BV�[�IC�b�e킎@�r����_E��3	�4<���T+ӗb��dC�T��Z+N9]�a��V�N*w��{u:�#�]�����FJ��-��/�ǧ_r2x�=O%4��r8����+�n�y݋��3�l�U.�:�9�؎�ş�eԋ����@�V���+ �Cϐ"ʂ�[R]�i_.��R�c'k6�����ճy����T$JbQC2����@�u�fjc��}�;��4;�)Z窨�� �&q.�ƃgJ��Ý�Co�~(���U���A?O��Y0BM� U��fʧ*�]�I�50G��u�e*�1$�YtR(|224�.І�.�6�c
L^��[�>���?��W��~�2�q�2pK�)f`o���cp�4ل�f)��D�eso��ON�z������c���r.z�7��rǽ�6���#�AwwoiO�d#����������<�i�.��\��\���W�7���V6ȏ�o����h<���B	r������淪������%A�Pp�%��K		����18�����0�0 �H�܉p�н��R��G��N�9��`;q�6��$jڻ������G
��]��GA�B�{�V��M���0�}3�&�m���;%;�G�Lw��W�յ��`�'�vL��1��������o�S�Hl�B��]Ӌ���_a}��H�/(�*����"B
�V��\p�����މ���e�%�&F���]�J�oK�n�V+���:�DbD�3}L�ſ�	#��z<�Џ��.X�au�yJ҆�}����7N���#�c�^�
:=-r��e��1/$P��_k���J/2���7ˁ���a�	-��Eú&L�����PT�{/ζ�U�wt�o,�YQB��v�K$����J-���9(�"ݯ6�5�f��a�]�&�6��K� ������t�v��-sI�{9>��AW�[����+x;nZ���R^+��bׄ�E�!]�>g�[u��()���mD �����za���i�N��P����v�V���B0hvAD�"V���V�S����E&2#���G��J3E��-���Zи�5n����џ	BDE9��­�+j��k�Q���L��n0�bg�f����I�޶B�rEO�w-��-�K�>��uS�0��@�4�/o��7 ��Tt9a�境ۣ�
CV7��E9�ҹʂXXDKa$+ �x3����~#0Y�w�jO�*�Z�{�q��_YV5��p�L��M�a@��ǈ� P����4"��:��T�T��x��G2��X�Ѡ�b͐�Z,9��[sty��OPh=�0�h��4p�D�Wg�]۳S� �=W̋��֭rMs�R������㕒:yC-�'� :K�{�g]����(8��	�I�ł�{���z՘%t��"���Z#��M렂̓�z#7���� T?�$�X�[��rrt�nhx�_}Ԇ�3�y
� �~zT��&�X����iYc�&ې`Vn/���*��q��>z/�!F�yI�i��:�}8��V�l�<҂'>%�0�C�õ����ޝ`��͜n�1O"D�����b[s���$u�����*"�0Ԯ�������-�s[�Ƅ��@�AfGw�-�o��Wow��BsN�mE"C���Àg���<��8�r��%��m(`D�g�=�7:>v��f�Wu�#H��VvP!�~BQ*\?y����%�Y�Ɉ��@ܟ�������o�E��E�=	�ML��Im�s�����i*r�z�Q�y�Ӛ��Df�1������4_��ɩs�D�V�b�Q�)��t럍�=���_(��5�^�n�Y�p�`8%mZ U���S<��;iɶ��n��^nl�����s�� ��k���%O�o#������eF[��K�22	������km_��.F��+A��Y]<L|�48���K'\~kwJ���0�;�$��J�8,B���q���[�&F	��e&�p˥v!�D�z�6���M�^۸I�� n]��&�؆��L�f7G��UU��<��ǿz��4W�t>[��5Ժ1��G}��f�=@���}Zd���6�1��0sΑ���7�ӹ�@l��r�+ڍ�*��E�0USN��ؘQO�q�1$�4j-l�h������)��Ԉ�"w�Wwƻ7R���?,?�s_K�%��� R!k�g�45e�s�I�$�'�'����S��i/��̟~�/�tz���F��R9qR��)�s�><���\���څɣ7�T

�;��y�����r���ȥe�F�?�>��g�	E�<�����4����}�.1+}}Mh���_KA�ȑ��󉂰�KA��ܤ�k+��ū\*o��0���Ĥ��p /�͓1��4&�?d���Rr	L��������͈�?�2�-ܨ���#�y�us:xh�����^9����*�b�UZN=M�2'�F;&�{��"�Z��KP�jl�ƿ.� ��gެ��c4����zHFce*�gm��ϻ���wS��$���z�x}p�v�K��a��V�s����0{�����2��
�>�x���6�5&`�AP�8%!��#�*��DQ��w:9���	��m�B���j�%#�C-�v�yDVE�f�����!s���'м;�j�p��ܒ�m��7�\^ë��u��~�:pq�EP/�����E q�f�-���!@��fֱC/X ���y�0�xU�tc�;�)�'VgT��U�M.�pz(4J)�|s���/)��3��I��+˦�uO���yE  ��Adɤ�iG���`�>�Kd>���1�K>s� &�Ji-.L�?q@0nS�&�g��ҷ;�t@��(��Dc�\�1䦲��+O��{�'䧶��Y�%��M&�U�9Ao�n^:k�.]��v���N�/&{���OK��G.p��S9�8�[��H�����i����/u��2�MZ9({��rK]	G6E���O"ȍ��,�=���n���&XR�G�P.�WS�#
+��.�Y^S ��oВ~}@�ٮ�n3 �I�������v@�S,]߉ �[��g�|+y9�γ��ئ��$�x@s���HQnX�s�!߾�b��b�5�Ll80�t<�mV���kFr]&?��JLRO(�~�6����M0�=�lS -%����`Ԝm.�̔��`�p��]ZWD�ET�n���o*2���J�����_ ��pP�w@!�7��:�%�_̗{����}�G��s)�HزS�`366��MQq�"{{��?�ES��i���z��]���O�^̦�������DD>��U�ǵ���*��<��+ḍ���"�	��Y��3z��$�E�I��Q%Nb�RjN]Ǹ~�%"�@Y�D �.-K7K��`�hl'����9�!���.���NY��Hm�Kňq�D#�sa�1B�П��c5	N47�*֦lK�i��YJ|��L�W��(j��#�B��b�%؈|�����kt��4��w�����x� �]�J0,�r+˾��+�o���Iڋ�v3���E�T:��835�	Q�PK�����^?@��I�xOK���f�3��x(�N�r(`�i�&g��vT���-�ƟO1O+��8U�H8H_�|������8ՙyӝ�s�p����c��Y�5�юdԾ�O�c,�K�v����=��)S3�9@H�l��~JĩV*o�dC?�Ze��K�z�,�Ĺ�.xf4�B5G�lԌ��1��gc&&�vo�^6,5�2�ۨ@r{���î�q��\��l�y�M̿F�	N5�ȖU�-�j?���Ț�����S���nb��tH3��J��a�.���B/b#~"�3����ژR6�Fq�6�x�W�(릶_$˻��R���F�s�1{)�m=�̥[��l�:�-MӴ��<��'6"�ٞYC���oR���"���D���	�F&�G}����E��Tr -bυ�)!>�,�ǟ�3�`��K�DU9�<�
�r�ň�Ag�G��()WU0���tAn��\`�+��y�:TH�l���L�cފ�1'�x|+���H��Ǫ�~���e��(�|�b0���3\o�U��s�0x���x�u�&y�]+��]�vV��T��5w�=N^s��Ǎ�E�k������	{$�nm�����dV��R��lRG/UI���>~Vug�{Iʷs�����|�F滞��[��y����ȿE�NfѾ��X��a�?��r��!D��iɧd�=􁗮��Fk"�b�Z{ �0�ESj��U3�Ooq0pOcb�U�c_G];�g�� o[���>���?Or\g}C�}�lbx�G�e� Iˮ���r!�����y���R��w�U�G
~�S{h-���4�w6N@��4�bi�w�Шj��֍h��d�x�{�����!��b���90a�%�0.��������&j��¡a�ZO�m��kONt5��m �R��=��2���ܺM��B��ݲo���<��Q���ɠ��\��Ŏ�~���N��}.����y;��C����O�d����fD�q�z;��f���^��:�^�JNBq���˗\2+p�%ya�[�;��pR�1_��6裣�eq;Q�s¦1�X����1�nb��7�(��o�rt�&'A◒�X���C��S{l�φ;�e��('m�	�](G�S����1��ь:�6iD�~Ń�D�ۀB�٪?��>l��2�a@�P!i[���o+�R��̓����+�����9R���	8L��'���lY��O��l�)��d;�"�t��ݭC�')�^c�uP��<>a�������R�vP�"ϝ%㨸�_Zd
=3�k�NY�J�����_��rpv8KKV�Y��J4��J1qT���vC�I����V���@��Gm��H���E�ݫTBȧ��^�����I�����
�3�[w��}>��C}�h� ��E�`����
$�g9�5�U�ү����M��8 ��9/���m�^X��Ȕ��������m]�Hi���LE�Ҵ&Q��瞒�C�Ǖ\E_8s�=�Ţ`��}?}*Q1� E�Ȱ���ͅQt�u}�*�xO���UC�{��>4>eFW5��6�JI�b.�}��rT���C	�`K�k$�f�5�i����uLս��N�sgtW�d��:OoA�T�AL<1��;M��tF������}͗��;nVqPIH��@�r���:�W�Sj�vM�G��T��'7�(�P難"[3�c�=Y=�w��w�X�$��_xH<�jJ�Z�؁��u��N��sҽc�.Ұ�B��1S�q�#:X�~�-|F���L�i�q%�$s;1|��Z�@W��^�L�T��7�Lr,���b��Q�c�r%�Dqyo�('w�\C��-�r�t�;�m�� �Oz/� ����P�lT��J�,�����S�#��3�]�[bH�;sY��0XO��H�/����Y*��_e��b��9�IT����&�l��/bp}�+6M�����:Ǣ/��FC��������h7��B��'�8�+u"9*
���/�_�@�^,K4#��p�<̐���0M�	�La���o!��%{��*��W�� �]�v��6(JR� <�U�`�w�#毁D�
_�rHuK�h�w�Y[	�����ܑ��^��܄<յ�O���	�����������jZ%��'[�p$����Lm��zwK��]�^Q���<*��Pw��WG���?~�u�k.E?�:��:fQ���/Ho%�#�Y��RL&�/�L%X��xS/�B����6{ѻФMH����<n�]4@�	\�U�c�!�pPy!���D�6Kj^C�(�Z�P�����z����P`��sk� <�e��X∵�*�|�'Ӓ�vE<�F�J��?���~����P���t�է�]���<��JLE���HA) 
$ \1Sb:��XV��f���K*�0��|a ���"���i�h���^t��L�~v�z�a���P��e��������B�`��a��u�͎I���J��B9�?E?�^�U5��hE�����\3��^(
ҷgի�=�閪&���t!3��`!u�h�/���P�ZTc���j"}!�r4!�
�v��I��$cB|gV�̺�U�aǬ7Ҵ�>� �dB&'fw� ���"����QU�G�p>S�`|i����T`?��"g�?��5���K��r���� ��#��4���ۇ�Q6�g�|�����2��sT�8�o�z���PQʾ�����d(���K����qP��	1r�����5��˭�W!�P�h����.�##��qS��ٍ��"��u`�~��Z�q��[���&!]�.�ڶ����ut$�%HEu��N6!�\g#S��;4B���i9t�����GZBW�]�Q=�N
���M�����v�\���j*�{�=Ƚv�SS�� nR+7l펰ӝ��K�){��|�Z���h/����o��e���
�����}���փه=o�5��Q�ݳYRu�s'	��;yU�=&������KQ���?l���~�iw{��o����7Pv��2ʥ� ��'�LA�Ⱦ3}|U�c!Q�;����:���i""�;��6e>���L[���$}Ouq���L�1�LY�d�1r~��Ȳqp|����%��c-a�@�rs�۾#ٮ��2�y㉈�/��?�~,H����@�cf� C�A�V��NE��X�?D�?��H�Hs�Z9��F���]��2�qط���U6	�g�4�/p�sM��q�'".&,��FOJ�b��8���� `�+X��
 Ď����R�bذ�v1ʢ��Cǆv�,3�SZ�8�ƥ�/Z �c�#�8�.�)����얍G�D��Y����t��7���J���uQ�g�Nn9����4�9sVd%�����������Kb�]<!�ȗ<C�@ԣ�V�ɹ7t$��q��&y�`c��������!�Z$�LG��+�n�\Ys�k�!�L�PW�.P��i&���N%���E��W4���̫,�?��*�D����(������6�@K}ܳ���j��G��*w�̫�HPWn��b���J���:*��=d��R����zCg<s�Px���)	�Ч�#X�*f9u��G��jv��B���!u8lFY�� ���w�Qkm��`��qP���ϝ�}yv�s�	x-DYYG���j$Ё�RY]
����V�:-ۄ�-�~J�2{AE�J� �@[k���)�7^^g��p����FN�S��~Hh��f�)u���64�m�v�r`��)+D��L@�nAXK��w򖝳#퀊~@��,��� }�Cu��d�� o'�3�2���:�E���"V��lT�p�Y�u�S|��)&0z{oS���z�@+��Z���I���&��J��-��"Y�uo#x�j�;d�z%���Θ�⃝�Q$��U"'ڬ~H0U�
��"�� @mIЍ�9(l;}@�I�6�u���Z��T\tF��Hf�N�
��+��H��X�{��`����ݳ���;d��P��R��	���?G�*���v�/��g�Di =�>%*"�+Ǐ�-ػ}�Aٵ�R�����(��j�I�Y"nã�U��Vwxg����q�p�ѿo��.~�6d�w��)>p"���?�ށ��23'
�vb0�%Bi�|uf�}I�̭�"�e�7�a6z�RDh+�⯷���Վl���~�ǩf�r��|��r5�s���j�~��w?̽�7�u$և^�������T�f���cp�  ��Y$�Tz�a�K��8��L��`S���Ŝ�ێ�R��k 3�"a��ӛt�ɦ�53�{�yl��&`4�0����l_�B�Jȧ=x�+��Md��@�>�&oh�Y�Q���v�{�ԏ�؎��@�JQbgr巰;�]������\Lj�A_�u>\-a�-�ŝ�.R���г�Q���Vv9�����ޡ�I��pq� GR����I�H���c��MMØ׆�#.O�r�U�@��F�v�x9����G��Z��S�П�>6���-k�_�W�Q�~�~�2�B�u{ڬu�����?�Y�Mtr�WB`0��Z�կ٩�t�hJM�=��Hӳa�܀Ҥa�o,Ϫ���c�:����j�z��<���W�,�ڬ|3��䒎ny��W�G�A:nu�!#��Z�1�r��|1��F�G�L���;�]��SΫHB��	O`���h�וn2/��o᮵����S*����Pa���Ŀ�u婀��g:�A��;�ak����'!
���+�!1;���0u}���f� ϶����w��¸C"�sњ�z�S7�,쿄�]_�P��[�G���͏�c�*��>:��`�2�?s�Xl�+��a[���⺾͆���;�V���জ�;�����ܪ3���/�_��8��8lŮx2����_���y��]���V���,#hd"�$j����g�-�r/��8�K�~�D���Q��y3��Ъ��㔄b�h<X�TwƐ�6b0`�Ӡ���z��2�l����0�ձ�N��%�{��:#0ު��K�5�7���ٍxݢ��>�;0��G�x#^�"��c�s���*�a4�⪵tt�)s��]��;5���DKג�2��֊knZ#���mٍ��%��e�1H���P��p��)] ����Ӭ����m�߽����ڣ�i�M�����i�myBm��,i��<��9_��\�I��վ������MKI�Z��<,T��`Pk.�ˌX��R��B�h�Ah`{��?D�I���؈��H�(E�o#& lϼ��f@Я��'��SCRX�UMe2�9�%y}h���qV�a�P�m��3J�%5CF�cP�:ŧw�\���g�3X��k�k!��b��&>?�Z�E�'�I���/��`<+��l�#��%ݹ�����0�_�p�� 
\?a1���2|V���]�V�Ã�+�?�^No�}G�w�r�C�nT %�k�3@1@!����c�4�xr���>�<?E�{��#���'	������h���ݽ��(��T�2�^�	 ��Uj�.��>By��9�;s�>�6E�EC�O�n�eAƓ\3�ks��˸n��wD����v����'VLx��)�Hu���[���%Z����}{�nl)���W�������	��
'�-�#�\*���s�q,ʈ)d�E����FP�L�晷S��*�XJ5!�~E�#cu9���-�sJ��wl�GO��'#c���ֻ�A+��o�S�T#��K	�˩�č����b��X�<��_%(��E���'��|mɀ�|nv{��c-tZkC�Q�g�����ڏ���+��d�8c<�և38
R�꾆.��l����؆��]^*w]{�k^��?��ܩ1�$�.�K,I:���}s�2㞊F�xh���Rp.�Q�q�^`ߕx�����(���r�A�S^DBL�#.l��7G���u�'�ی�Ќ��a�����.��`�$
��x!6M��\T?a�(���'85Ո[l�gY��N�i��N�����y/y[K�r�H�"$�\D�ɕ˛��v7�-�u8韓���Q�q5/�W75�m�(�9��>�c�n�賳�U�t#��[̑�xH��{�Lv(��#@��ʎ�B99��痸�D!L5h�xT��ѐ��r�d^p`���6T-�l=�E侀�A�3J�Z������[�d���Uyfhzo	�(^�3��^����X�Q��>>�37�a}�|��9�\�2��Yc/*�9!B�?l`�)趣L��C7G?ߌ���n��� l"� _��翿���%=S����6t������^����t�<#��eHG���P7�T9o��YH�*��|�*��g5�u���%�Q���4ɒ�?/ᗊ�y�a�y������'L�V�!�F����x�0p�6=2�����Mk^K~�̸��A�Z����ӹ���s\����9n���b횧������oy��d ���eNO��Y��G�y��d�W�B>��q߮��;�Fog�����^��r�dl0���s_(ƁI���D��ܣ^J�F�0�Ť�b���>*��({������g�`G)D����T���K�$*;*��C0U�Krz��G>��`w��*��"�CxJ)#������#�;Ox��|똪�z!ϱ��4^�uJ�?!���;���)�M��Qv`�Z�`��Ā�E�Gc4�ЃY���7Z&;��?�&����D�(�EXx2<\��L���*�l�["�<=B���+�۫_�]�4q��/۝�w>~��E�I>_4ԇX�}R�ό#���oU���g��&b_1`����Ǌ]����~h�*�Q���M��'���	$���䁢`)Lsz����'����#��C܋�R�R����=�)|w����G�)̸�/P���E�4��|%��Z��0L�w�j��,�=sz?������S�.����L!3�獢�p���e��)��'T�-�g&�*XG�0� �iT�Ao_G!�l:'��:Wl@*⏗9i��P�Ў��L��V���9�)S��!�_�0/^xz&�9?B�������i��J������зbd?����	�A�0X�z��cc�?�j�P�����[�}}�	|�n�/A�L��n6��?̯�û�_Ē}��1εY���}=x���L_.�P�at�m6�U��)��Ih�a��o s���;��bmh^���;�6@��V<g��6톺�,F�EuN;�~R0<�p��v�ަ�W��������u.l�ƾ�L>xO�	�����:��uT:���֚N) �ND�&R����e�G���$���z:tP��$�e���_uÞkxA�ʘ��C릉�� ���
eR!]�Ի	 �[jˏ�T��̾����g�;Gjq�C	PE�%�tt��1U���Y�ҟ�bkߏ���4BZ�oi��vz���d��x��$�Ko
Vk����SQ���i�Gn���K�b*���&㮳���]�j	~h̒���3�5����7^Wm��ssVܟj�m�ң�Ũ�)�;Kk��A��Hu�6YW�-�|v����T�����j��:���KѶ�Ǝ
$�2�yG0�T���(�=Gh�':.��M���·`�V��X���V]s�7O�q��f�/ AQ�~S|.��p�"	�8���� �,�|��z\i2k�f"�I�!��|n4�J�`������2��\��,�Hw�b؈Rd����?��S���/E�1�4U�?m��Z�=��*7xV��.D��I6Qd�DcI�:%��'e,�������(���$����҄�ϭ�
n֨ƇWxl��0\NZ�/�2�ޥ�ν5���V���s�5Ȫ�r^�Fz�>lf�1q�����t*���S�������L�N��1��	���7�B=�Bj�NvĠ�%�]-�a��c���U�4�ی=��ߴ�!Ŋ�7<����r�'�����8B��<N��I��D,d �*D!��[�g:�����_��9`�W���r���㏳�������RլS����{;T��dȖ�DK��d��%���b�����z��T�j�?W�@����Y,J�JYd���É��?�&�lu	`����fm'c�T�f&5��퉼��&���Hg��5��}��)e:�Z���Od�+ztc�Yq#|iz���7��	�V6�aǳ��Y �m�i�)���$�����`(x���x1_ުx\����'�S/&��_��:'�4^塋�I�g��nG��N{�C�98sk=\�z$���fi>�G�\���H�b��C�!w�N�|����-��������X�Y�H���^c		��?�a��?�)~�&,�	�T4���Ѥ�L�8�\YG�ҏ�Is���F��[�"��u���,�f����$�"�?�s^���݅��4�>	������/c�;���u2�^���)9�]�dA"��vT�K�7�= DZ� ~,����TYyY�Ӊy<����I�H�[�xY�5�+VJ���֠�Ԡ!/崄� ��8��"��E+ez}!���Vs-���n}׫�Q@f���@��`���`N�	0 N�?��+0��s�~k��G2BS&`Bl�dy#��]a�6�{�����i޼�><2�u�p���	D�l�B�͔�I��>���tZ�wC��c�o���_Z;�s��|�I���j�M��}\��V0�{�r�G`,8�L��L�Y�10;�����&�'�H���'��ZqٙQ�፷�+��s�Tu���j�ox����[d��/�$��k_J�+���&y�>>��s<p���!������Z��u2d`�y��h�.�NB�S�d�W<?#�&��^�$��"��ya�@g���2 �#{��9g�vD�۟����UE�s��q�Wݪ�
�;�4j�2��1c��ko��箞:iw0,�H����4r�c�`���a�8Xn|����F�Z�p�k��������T��׮Vh۲�E�A-�����Q�3�q��~3�A�^Q;�ӷ7�q�|O�e!��hXlx��9w)��16��h�o����/��{�H�[�͂ӣp�Exl��2�����U(�4f��o`���.�i��y���tW\"j	��~%_F�4���,u�a]G��e$A/7�C�lڀ���y�c��D���*�7@F��*�b��9Qy�'H��'�=l���1b���	���T���_�
n��>B�A�)�xO��i��4�+����M���`��8�^��7�F>
��R���l��ePHZM��8��LJ��;@%��f��6�����Ǭ��a���L@�����13.u~KM�|gMZp�Ky��\�6+�b8�~X����+���h�w)��.�����ʻ�h6�:�w!/9
	�#���. ���.��)�97�?%�f'�k���z_�j��"!;�k�X{1Ig�R��>U&�ҚS�zSk�������*�����F>��h�,4�VO���Ѹ�<���{���Χ���4��`�%� F͙(|���>�Q������I�`���o<�{v�d����/���t���)������E�%�f�ݑ�f�'��zlq�'���@«��_�pM�|	N��S��%��%B���-O��1������4)�L� )��bJ�?����8$1k��ǣ_�N������l�t�?4�]q\�5�Xv���G7|�3�6����e��7���u��G����i��Zx[����Z��!�!��[�����S-�}p�u��f�ؙ{�qLQs� ���Ԧ���o8kOcc��% � ~|�*~�E;�}����d�ɭ��H���Ƀ�=�J�Z�s;���4�7��Yz��Z�����P���]ĕ�%n���]ې
�m`��pH4�����R�8��!Jh�{C���<Q�&m�A3����*g��U,�X���������."u�r��\�I`G�z��BC@ʏp��^ڢ<�c��I��2�q�8/�Fp�Q����j���7����c���B��/3P):h�� �LᕎH��3W�jfO�wc<T��6�����E������]d����z�R��#�i�0Z-�8���r�0�
�qƋ�,re[WP
��Yb��2-���E��^��6>�S"�S��~�s�(�q��{sU�����^�S�]�� Z���BA��+��A0h�j'T6��y����/d���iJU�;��"]��_���� �6F4u}�^/��˅�/,���կ��E|m�?L>��U�*��D*C�K_���l	5ښK���T����ӕI��[0D�v��W7l�.Ry��L��g��SF�������Uܾ:U��'��``��]"��/�c#f���O�V�,)����G�Ka����;�M�&jL�l�sZ\�L�������@ ���>���o��B��l��Dl�(�v��?�ڔHFT+����.��� ���ư�钠��j����q�W���B$$������'���#��o̎?�w[����݃Z0мb�ҍyL��?)T/�il�������{���M��4�Ot^]mow�
{�lGH=��}:��蔙�=�A�{B���Bz����Ʀ2
�s�v�w�Q�Goa��E�-�*۔��5����1���n����l^× ���H�7���㦝b�J�p������3��v^��"&v���V� ������3ip��W�8�˧k��b�m�kc��4����3�^�#�����qv�3�j����j	`8�*HI�냝�Wν)3)����-��%9u����w��PNޏ8���������I��cD',�?�ۓ�<ñ��ZR_�C��w
���2�x�ހ�bj��p�$�i���^}9�Դ�Lb
�h��� �.ǅyǠJ��� �V�(s��f� lfY�oN&������>r�.O�t$;2�Ô�Z���\���< ����͝\4���*A{�� t+��{�˱��Jw%�4ͧ� 8��	l�l�dB��y ��.l�{�S��{����K眐�ۂ2A��n]�U�8�r��=��{[�#�Dg������Qy��>W�;:}��ӷ�d���S����,_M9��9/ی ؝�f1�#��n(��1��ZZ`�P=t�+͇�adb|�j%��=<�*�z��#��==\��	����`&t�;��+��z:�2A�2�h�ye�)`bY�%�Y^�������I���N�\C ���L��z �]H"pqP���d��֪��Rn�?Y�<�0E��������� j���$�MJ.8aʂ�Q�Vʟ� ��m��.l��c�ot8[�NM�=촱��!�$\���g��殬z2�(�1|j�{�R���% r��f�i|��	����D����7�Gh����O��r�B��6OIS����C�#�&@U��k�Q��P�3W�׵'�FE㵊DB�Q�lG�1�6��q�������Z���8�e�?z��\��B�Dn����dL�]�Pa�E�x�&�"-�L�Ɏ���䈘������5� ���Ҍ��c������k�+#9�/�jg�}B�18|��z������tbq���\����切-!&�έ��qKY��=q�&	=�r��E�;^�,v�͒��-�)s�E�Qy�8�a�1���G\F�Pܸ�X�%�>T�mO�J�Qze�`�z�>A�E�t ^�v��e����Mc0�RG�+�4TK���*LF�o�l�\g��KR��݅9�y�fxGA�pTy:Cø`K�8#�_P�'Z��6o�n"���g�!���y&�b��V]����0g0�}7	�:Ud�`���L�dC��c�7��sPf<N�P��MD��S<�����5�j�3�OdF
l�6N���=v�F��nH�QYq�5D@��O�Kz�X�E˹̼�m�KB�h�K�K�_��:�
іҜ|�n�Zj�%�\�ґ��hl�r��^��'&� ��v@G~Zdӂ|���]�J��W����j�ZzY.l�]�K�b��$���bq/�ʕ�n`�(�O�'�@�Y�D�*h<Y.���e�ed�A�u��j�佃�
��{�FwS1I/Ėx��j��~�!½/6�ä9�za��!����y��T<t71Lf���9��6j�4��V��Z� M��SH�`B����槲⃰��] �Bڳ�_XS�Ym{ѽ{��hn��I�
_ }���DG9����X���smr,s9,IN�O��Wv�A�K)���c%����0�Tl����H�a}�C�e�H�����ͽk�f�J]c��L[(�3%��`/D�>�~��!9�1?|��}D}�h) ���atR���זr�%��3��~yS��"|YF���qy�1]�+pg�lG��i?	�LG���e���p��D@���v�&�2�ﵹz���%�>���`qc{	�QR�I�x��\ϑ�#!�x\�gUk
��3�5��ǫ1���L��(~i+G���C��c��{��/�_�*_� =�8�/�pT/X{��̈7T��9Wj~׹�����`_�b�����_5vZ�T����K��̓6'�鯙�/k�a�����ᷠ왼~n�o���!-�m��Z���X�_�й�BY�TR��I� �C?!BqB?�����`_���ϒ�C
�fld]��Q!�1�����E@#��ru�WMz�w��Y�( wAF�St�Έ�m�Z�S��-]>��E��P��\�z�@I4ƠA���k���x~z�?͐��un8-r;s&Ƀ�x��K��XE��_gbSm��}Pwo�)�(\���w>�������4cj٩���&��/��a�ó��q[��_�x'�� <����59/uYm�(9^1Ԅy�
%�M4�O�����N�]Z���Z�Q�i����OR���r���M���VD)1<Į�Ƿ,���3�)�I�~'� �*E�<�]��E��~v/���ƭ���Qإ��p�3��H�������#��h��7O~+�$���1e$�KY��z��ʳ\3�m=��RXx�az�p�����I��s���ރ�E����"4��
�X��c�|�s�7��ą�fJ>��}E� ��D_}w�#�&�tߗ�[�ɣAX�~2�Q� �k�$�4��"��^�%��Xc�]\��X��}�n*��3sٔO&�ԡ�����o3�&��:�4�ddU�Jgt��1)����{fFu�1���e�e��������Z$;)�szC:��{����ɖeZ�ݜ?i�X��Ri>F����y�<F�˱i�aCG餶�p�����=k��z!������RspoLf��0/���8]�)uR�~v�ʤݾ7�eϨ�㓨0,J�ס0��?-�a^��?�R�`_��p�2ߗ�5|6T8d�r�_�EMr��.�q��4�u.�$� L�����w��.�ɣx4�J]�]W�_p�[d�=�ԣ���]ߌɂ�-B�t��=\`�S�\��N��0��Z
���9'�2��rZ�*#y��V4JW����߲��_�M�� �Π�&����~]+��6�߼T����_{*���h���C�~F�5j_>s�:�-#���08�*�.�!���t�g���z�OF��c����FߓI�z|���:L_��;^x��N�L��,�"	-�)��e%�K	j�`�*�����O8��Y��AP���>�)OC��'�{'ˢ��G���z�U�2��+q��(%�+�D� ��z5g��*ކ����o7��@��%5 ã\o+6�+�`萌��41bB\�}���%�%����~2!�>w�$�w:�,�'� ���Ƭ�]��]e��];��欏����
뤻 �ή��4�}���pɧ��&[��p�k�BO~�TQrJ4���5P�b  F� ����K�
�^�C<!��ߏRT)��#/�|P�������6�Sj�g7 �Ђs���������Jo'���E}G�jؾu�_���в�����.�ȩFxT⡒�M��ݔz�~Ɔ\�$���J逕��� K�9��m���4����/��R�`�T�N�i�2J��ш���Z�!���|��9��g5�[�zl�1�/��`ˑjq/��y��"C�2#��FD����f ,:�/��x���H�nr�CZ���xݦ+��xQ��Jz��XR��0��>V�i�r �f�'���,p)��B��ω'y�&-HN�����)���٫M�����S	���h'��:Ǎ,7�N�!�`����D��K��set�P�jo|�wWL��Ж�b�BT���B��Y/њ{u��6z����&D󨄲��:��T��u�J��z�$�EM>2(S����.�3�hF����ҝ�)�t���U��tN�?�Hr���D4t;����-L�ʅ��N#�$������#��85��G�y��ӼLC�kqJ�d1Q���Ke3�M�£��M����b\k�&�h/��9%bj&��A+Պ$9�'H����:�-P"�^�~j��� �4���&���=e=W3O�����c����Z�9��Z3���'���3���rK�(in�o0+g2����K���=ꈷ��0C�g�o�|L�c��/DF�_�Q�:ӣ��t~�0Ґ��"�;x|��u�%�Ԁ´ ZÓ�4��Y���?��:Pk�4�ܮ��R��ٽ��w}'�7�k�{��
.�.8����-��4��m-FQ�.�>7Z82��|����4ǘ�|� ��7�TPȂ��}Ӿ�Į;��� �uX�ES���>���S�q�g��~��	�3E`�킱���aT�K�oP�B�w=�#��:v����T���̣������E�=���R��L�zr��h�.*����n���[�-�b"��	�Y{� �`�"/�7C�{!CG@3�����s�P��~@���I"R���2�M�~r�q�9\����O,w)�Λ8�?+l_���2�(�r���6v��c�Y�&�#�raFg�Զ*ݐyVo��".�&����GG#�N���b*?R��*�A�{a�
�!�Bd�5V�w�B���,b�p�Ne.��_St '�|��膝�}9��P�:���O�y<* ���� ���h@~��O	̼��ᐌ%}��6��:B�9���x{��+iwߗNz;�r^p0�ۺb��f0=�������X�r�3[ɡ��vVGLd\J�Q��u� CJ��1m׫�p87��BXp�O��pPsG���7��IOdG|~ ٯ��S���'����J����O�t�%9	��t�AwJ��𹡛j5���\/yz������b �ec�������&R��m�@ɨ�7"gHOFK��Dݱ�Z�K̵N9N���J<���º�XbP(rY���¤�EYHE\�I8�EWkR�$f(i���p	3�Z�h��<-s�7�_*�U�X���#w�Ņ�u�\�
Dm൚��r���h��2�P(͟f}q�1y͙��*����o
y[���*^Gr�NRP���Ib� ,�n>�z�:�C�ju�b;���D��C�~�@	D_覉�W�2NfG���?�=଴����G������������_�7��J1w����P�h��t0�3ѿ�D�uԶ�D�"!�5��2���&���;r/s�46l��.�=*��kL$��f`��L??m3>�d�|@��Y�.�V��i�G�>�`�R��H-�lT���	�C%B�!�đ��>�/}�b)$3&���r��\�w�	��e�ؽh���!�����E�X��9߳��1�6=u���C�n���+���!�a����#�>�c���|?���xʦˡ���|X)�~M���O~W�	D�v��_�^_t��C���kd��(�ܳz������	~�}���*���=��ʝ���|"@�R �O��n��×�r`�~�D��~L�mU�P��f0��v_�S�L���p�}L��A]Ws���JEm\3Q̲��(����ah�Ӫ�Yn�������~��`'QBS�@�c�8U8qM9Y4	�Z]���$t��[�I����G@��W�{\�%��SvK���~DT*�>��ڊ1�Y
���ۯ��������P��Y
Ł����Ѵ�7<��!�1��"��sO�1�~�p�h���u-k��]I]-����o�z�!��J���HBT�Ī��ש���$�,a�F4��d6wX�����M���\���״,�q���u��9./��n3���?V.��1ҕ~��s�����	����%ޒ��3,�s
���N�d7���]���Y�I�u�'V/���J�j�̨��b,���MF�v1�!������~i6W��;�>�@�▋��ڐj��鯴�;>AH8E�Y�Nlz|q�n��q�菰qh]m��;���S��DGH��}�!�D1x㟕�Y�3��	�Q�c:a%;����H��"����+X�q EIR��l����#uh�YZF�	�࠲c�G�� �5m�H�b�h���|NTE`+��������>��Z(�f����b���?ː`�N<�L�E��
�Ky�e�>���'*��`rY6vM�yZ�a���LZ���wb#�{]���8m��'�Pl;����iE�Q�Ȱ˖4�1�w�gvawc.f#\2p�X5�?*d5��FQػ������UwI���|�AZ��1@�p���
��?��`5(�*�:|�_[�F�o�RE���,4�ʠ��6�!2�[�����Δq��#��l[ū$n������r\���<�a;��kT�����=�oYCg��6闥}}np~���R���p���#�� �~���e�ڄ�v=׶��+��[�V��r�_�$�F���/澨H�>�P\-tyB�_�M�h�١��S���\���έ+ޔ�=�&X�f+r�@@��}�v������{��22�XS��罊�>����)A� Aϧk�u�����M	�R�j���4�$�ޟ)�mwyao�����Y�n�}<�{N����52���=��o!&7�i�ߎ`+���q�w�8
�����U��:@K����SQI��4���a��D��C����t)�tM��:W�z6�����)�)z���)�*nZ+ģ�cl$�qI1Z/ '�H�y9�}�~��M����.��a�,d��X/������vL��T�g��������LE�a��3o����;������}�S	1�lV��ppa��cH������[�h���eJU&]��}K��1�@K��z_����@�N��K����&�
�g�\��p�jC���*�A�I#%�Y�g%�#�s��f��}m8�ɟ
�W\�� N^�l�5�w�E����V�J�|��������RR��Y���T��c0n�{�g���j�vel���ϝ�|�NN�C�W��Q��؏��YU� U�aD`^G=��m����	=�\P8*Y �u2��VTh�-����Ŋ��8��_��5<L��eE��ͬ�|���g�u��tĪ��,vU�vy�O#R2�JLy|[�4`.�f�|e��aw�/\�7��x˗�)�1�<��E��w�`�4b �<��w^J1B$�#�&s?��%A���@`ɨ���>Lk����
˲��\�P<�Wo�!O�P
�PP��4�k�yş�$d#���b$c��D����s�)g#��ڡ��"D�K�٧�s}9m�A*d"��tFBF�e��x��JB,�>HO�]��*���?Y��I����O�h>��������,�H<��)F��;ߋ�	����������z�?�<������-�@��X���!�tZrbZ�g��!��/���C�{��Kص1�b���X�������×��~"A�,��ͣ�~�K7��g S9�j�,����iNv*�� ��,wB�7
 �B�p��_��R�������^r}���V�h4�,<�ٌ�Is&�)���m���^����T�]��.!��-Ri�����	Iie��Vu��%�  ��j���t1��w�pF��Wa��C�dsu*��\������(�H:d.@�P�����I��&�Tu�?I9&�ů^0���4znUj���Gۯ V��~f�n0�ɂ��MO+�<_�b�l�݋a��j]OQ+�(�(��t�g�F�H������[4����<���cm,2�Ŀ; ����z�'��K�%��+?�`^��j/�Q�*��gK#�k�I�C��/j{v12�	6gr�4������1�}�y�x
|~���e�F*e.�$=�)ħ��O]�������c�Z3���7�K)��hA.�n���X�OQ�7/�ô��L�S����z���4���4�����X�z5�ց�	>�!:�1Ʈ�����۔�����gV�M�s����d�iB��~#��P���KΡ�äCEE&U�KmnZlZ�H1ijC�D�C�����"��Q��DeUM�J5�}��/�����i�[BK뗙�<ն�8��ۭ�+���տAo�ͺ�k��0	�5KV����s5 ��`�g�F���Kcܵ>̀�0xN�=����ل��V)�^o]�L���0Ҕ����qm3��p�D����`�88"��'�C�c_��n��-*4�5��7��&��T�n\�����.����)��Yo	��ID�E��:~8w'W��2�-��� �'���ވB�q�3�8�Vw�F_)�y�&�?ğ��:�1�߇R��&�Ut �7ls��V��v���ʯ�[mC_bQ�����=��c]��	�%���a�&�md�v O5�DKId���`�w||�mb6j1�h���Td����:w�����'
�<N����[?��WׂU-$-��D�ʖ?���Rƻ�1r@������4G?\~���Ux͘���R���5x�����*��Zt��t���>[;�w2�7�a�>�q�fhtՁ����,]��s�Y� �%�l`����@)��Vn�d���D/�Hb�0�`�����lz	������i�B&֘t��Y�#����q{����2CR]$�bs,��������[Ȏ%s�� ��,� p�G�u ec/ωK}�%ؒ�N�p����~Ju�\Є�M������&S�j��ʁׅ�N�����p!tP�o�+Ua������~i�J��<�/�x&�;TB�2OC���p*����(�!��;�$s�*\PR��%�
]A'��4?����N]F����]��b�/CA&���n���ʩ@tȽ��˧̹T�ѷ~c��.�%P:��ű`+�'�5��"��8�И��}$ c�F��81@�/VZS��Q�5�QGqO�s�=Em�G�]���<*���5�=_
-"Ѥ%�+}�v=�����51s�%���P�1�8O���I%�~��k�%�慯o�oa��{/`�i�}	���u|��dv�9����.T�%d��>s����^���s�Rz��O�7�,�*�{3��U�rb�NJ����osyDܟ5�и�=MB�ab�IX?����Y�\mam���"�� ��9��o��h����<p�3y�
J;b^J)���u�I��c����`h�P�?���r4b"�z�l�w��@��<U�s������Yi�O��!�"�������2�A�zh8D�_�$�,�J���,[��.�{;m�J���@N�+�}](B�~�}cvC:�)�%��r��O���ꇥw[U�*8U������O@x/�?�"�u���rV���h2���2/l$�h	�&�ۉ�2Ϥ,+C­up�Æ�<k m����n�إ-��3C�({z�5�n���[�'�u�x�
(��oKn���7���o,���a�B�>J��<���v�f�����N���9�uՕ�mv�f/i�u/T ��m�to��2�bυ�6C# �˂�=���l-_(LJ~jbri�-c�="��9�g�c���^MZ�Oz���Y *M�B�Y5}��l؃j�r�~�Aq?�?��c��D��RG��2���v�.�w;�A�C�(��&�p1�~C���6��ip�%fa�n}P.oGZ����.�+��8���%�Hl[�R���T�>�(*˥<oۊ�ϓS�g�u�.s���B�Z��n�<��`���V�ލ_r��M�ͪ\H�n�O�W���X6���{��[Yı�e�8;(f��٩�x�GiT�ļ �χ��jZ���ؔͶb��1�om}�L��oZ�g�:$��P��<Xp�@��:�����@�~���j||�A߰#� ��A&:�
 U�z1��c:^�]+��kn��LI$	o��uKxCu�����㷫ej^�:k�.8������\q��KК	�/}e�>��F���{��NK��a�Ud��OF�VYcY[l�գH{Ah9�� ��2��X�P�W���{�OB.�'��ؓ���S�Y�n�J��2��N����?��I��GOeņ�9�5��9�>���F4�Tq��������$��V�hw+M�Ug
��a��RPׯ?���L�l�' �}2��*eI��g-�5�ZQN_0��W&�`>�X+]*�L�9y��I�Q�	Kq��V�(�,�`�������z%���ag@D���1�����	mT� �}:�'��a�,,Qܮ��s���'q��Q�_k���9 �6a�C�q2�����V\�2�ա��8������y�@qU�Ȱ�d�~��^u��;����?��}v~V(u�����~kij����/Mf9�79]��tCw<[/�n&EO܌t������	C.w�����hz�d���k*eȪ9쫤��E��ŉB����Xe���RX)˓I&$�ƺ�-$���!���vk�y�q(�tX��׬�B�'�hF�u��KI�l���l�}�U��]�T��l�R9k/��.��Ԗ�^��E�l�+]�xk�tp�7 �)L��6����߅�K��e�ш͠�aL����/�|���Bp�Wl��ڕ����K6τJq��B��H�E*p���z�֥�f�֑���5<*͚�ʫBW�M�+�@s5���R��ѯ��,0ԩ�۹K	�; ����r�Ѯd5N��s�Nw��ep�F��'��}gc�Z6=���=�m)�:,p�.����Af�7Q��8O5���)�$�,;v��in��T��|�d;��X����9y�-�!�0%��#�(z�����K \��~;�` ��I��١�$�ݤ����OV��4p��
ͨ�(�����w,>�\"À!N�i��}�h����b��c����ޒ�5�<�_|�	$�v���6T�&��d�2*b�d������
��|=�,�E�AgGu¤r��&���u����ƚ����iϨ
|�aE8"���%����^���(��=���
(RҨ�� x�3'�nlȆ|�i��
!)$���U��*�#f��)�G:�	O�)U�h%!�>�ԑ��{���,�^5П�Fƣh�0�2�a�N����p��(�2��I�:�z|�P��+��=R+X)b0c#�w�L�Di0��W^z)̻�J���-�{k�^(I\D"F��D5���\N~F�?jXD��-ƛ��?�Ǎ��ۼ
P2����:޶�uRO79 /��0:�%T3k�	ei����Bm2T;M�,�[�����Q��$(%����<c$�� #���b� �w���ԩ0l���W2ۧ�yηL�������0U�Ay�5�J��sM�*z=�^w���Z����Ǔ�oD:[l�U���O�'h�����DJNtee�d��ZT�N�ߵ���rp�����0���ՀK0��k|�H��+%�6!L�?�r��1w���~�ͧt�C���*~RYc�?�O�����v��]�ڊA2����y6�ep�0�pWsf�'�X�Y���w5��T�L}��}�u�=�32�4*o�^�Y�1ͷ�Mݬ0�#�����4_su9�9�O�f�Y-o���~��VҪ�j�C�r���Bg���ЪEA��Y���l�Q�������V�yA:�ϲ�`�y��4�P����6!^μW��y��ᶈ����Dq��t�΅j7+L�wU��=� ��l%�2E��	�������7Ĵ,�RZ�3!V��#�����'����]	V*�&�9��n���ٕ�z����R؊�7��$봖���n���o&2�,h�fq�:%u�W�9}z� �2+I�<>g������P�N@���c�%N����\g ��]��ɾ>�ɻ���VR�a���*0Ǝ�����l�/��i���Q*T�G��m���C�?b]*쮶-������H:���b�L�
����xw.L6w�C��?c�ԼP$ЪT����(~�ͷ�W,g��I���t�V���3��M[D���i~��5t����K���i�O �پ�9Zџ�Wp�f�Ǜ�d,C�"�h����X��f�ѹ/�c8X-����l�S?�� H�t�<�?h�BUI� ������U��}��=j	C�lq 9��蘃�S�5�j�#p|L������Y黼BV���ԛ^�l���X�y��[����A)�\o '=G<5��z�\��Q��=G����R��������KG[�E�mQ#!av��y��1���$�<ϳ�W�`~wV#��w�����Tf�*�5��}M�߯<+8N8Gt��#SZ���!��ns�Z����;N[5*c���?HoO�p?��gմ�`j�t�ݢp��Ǉ)6b�6I#�Z�����j�ݩ��ʤi`BRC!�n'��p�zjP�֮�P��K�&'��r���>�;�����I�n�
�����R�jº����H&���$���x7'�܌?w]�ohf�BѼ�!�u�Զn/(�`�."w+ʁ�$��)�e�G�ig+S�4�U�^Lg�b��Cз��W�
Q9�pߏ2Cw�w���@���F"D���U���pY��.-�G�F���n�����|�QK�>;΀�kQah��U��8g���"+����vA���s�T~�#g}pI���
��_!v�=��U�0�����lQ�+b��rBH��P%m����)���������VV�M�r����0�T%�ӝ��tR�mb�R��⠚�%e�-/�T�lN +�Y������pn�Y��<���:ĺ�3��xx �`�g�Zxd�����ؿ}ϧN�,�'�%���GS`���h6K���/��/W�׮�Wx1�Uq� �;V"��'�p|@�5OQ:��޼4A�ĝ��5��6q����x>��6�.����^��%���qnj�:�F�ɳg\	��FL��t�r�A�5ݜ��D�Qѻe�Hَ�I_H�Z���Κ���௼�^�}�Jˏ]�j���8L�TŐ�g߮�����vߘG�?�-kb%��w�CGZ�RX�Æd|���NS4��� �P�ǆw��zpb�YX/��į��\>ˉ�eǺ���a3�O�Ef�F�בP�=ѻ{NR���@n������9��wf����b�4�g
��*�U��uc����7�5�ٟ�xޞ����1�w+Y)T,�fK_�`S�����z��æW^�Iʖ�/�'�$fH�˙��Qߥn!��>2-�/�1x!r/R�g���'`?�NH�5�b`
(�(��p����qȴ��>13�Hdv�����#m4|h�}�@!�I~K����|8���}5 p���Hֿ�����׊��X�X!qc�a��|ؖ���w����o���C��ڝɁ�f<֍p��0_F������1�0�ܥg�%pū����/���.d0�����f�i]S�g�i��}k�r��ό���������]K�G�A����U���W��ඵ�c/'�	�;�<}�P�F��^?�)��ru�3�\3��%~��;~��OEq{�����HD�m�~{.~� <�� �o(��z+��\d��F"e�O�Â�Q�=���=������/�D[A�/�3=	&ɏ~��>��C��!k.:�;q��O��IyD>v���Y��F^��lD7����J9
�ǥ���Kp[�с;RQT������If�UO��`���v	�X�/#��3M�|������{-J�`����<�EV����[�_��&��O�z�������Q`��T��-¿r�[T�+ݗҚ2��p4��[�عў���u�2dl2�NŷKAb\HM��ǋ���i�)��%k�τx�������.Cʴ�����U�c�����c���d���I44�B��fH�u"k6��oY��!l�t���Z@�=��c�P�����֟�(��}�1Ȝ�ߪ1I���д��L]�'��	R`*�)O~r-��;`V�&c�ߟ��S��|"��~�\��ѣ+c�V���+Ɩ������t}��=`}��BQ�8�!�=��u�ۮ`IOfb;��]�7eNW/zu� b~�D��|�����+�W�Mu��6е���O�����-�=�6�Jg�y��o������ǞJ$Y_�z�0(��י��_�#�`5!V�UӘ�&ߜ(@!��	��0��`@B��4?�-v��6Y
�Pw�ͩn�Yψ�+y&B�d���F�?��SM�f���$)��+�Zu4�G���]�J5M�GUT��+���Z���v��j!z��E�]�x�xG��5"I3�]@�}��%n�\�KNR������U�i5�Y�Y�R4#W�ɘ�|0��u J3����$?aZ!qS�D���k��;��1��	��a�K?d+�҉�t,���A�~{g<�I� ��G�l��,ةڶb�-4��*La9�1��3x2ai��Tc{�삹F�������.��6�qz���s�e��|S�,J�
׽��U%^�B�if$]� i�g��B�:�U�����	���P*����P���7͍��J�N�LYI&F>bYw�G[}�3�'){����["�i���)v}lLM���$�p��S�����
��_U\�+�� 7/RsȔq�5Mϊ�Y
y�/h�T?���@�8��}�O�إ9�/��a�_��V{�QUQ��'��1�JA��������^�k�S��I3���G�M���C0�1�y>����}񧻦L!JT<��X��oi�ߚ<�B�B����>d�oP�����K�ѓX<	���UHEP��/vE��{�Ă�$����V[�}k�b�����w���k@��k�>�ng�F�=���P��S'�����'�g^����\�p��#3���t#�-�����#f-( ���cB:�v��G��!�M<�|l[�9��w�"��	ʺ��Q�)�s�k����T��6�z)'.�U[�VDD]ѥ���qeS\ ͉U�*��@��<_��ƒ'4⛳a�׬��b��J�p����(���T _������w��%������I���?����8yn�A`��,��{��b}�z��j,j�C1��"��)A0�v�Q�����1�M����!8��Z������#�<+O�t�����K�Q��[z\�ژ&��+J7��$�=\�jvᨑ/J�cY�O�N���mnh�⭼��I��İ8i~	-�M���qܗW#G�:02����F��ͳw� ��-�'��[�5������z�?�dY�������|��5�3�� 9X�e�k"��}�M��	,g�E��!��\x���B�����_�ˮ�ؾ�^���������܏�F)bCl�w#&��Ĺ,�A��G�Ɖ�@J&��3[�0n�u�	
0D���iscI�VD��g�
qo������\_rH��ķ����Nt��OqFa��z��"h�kV���OH��9��,tŻ�����bbn{�Lm'�1�Vf��)�]6�"�<�v���Ud$�Y�)��ڐg��l�0n��g�l	�Ts�s���(D�8�cH��E��U���*ԯ��,��>0�z!Y�O���sC<L?��	rbЃ5�}>���b�?xm�/��B���;B�O���j�a;N%fsi���0�R��u�ΩZS��l2�M�"�`�7d�y9j)���&�F6��L�Cr=WRM�h��m1��/^����`:+_�_J1�5����@i���3%�[x�B�5L7����}�A�j�Ǔ�6�������*� �}����ߙ�.�ڿ��\�A����O]�����]K����B܏���8�3�E`�t�7�U��Z6��X�4T��]r[Z�	��6�p��O�,�p��zߥrH�8T�ݻ����E��6�и���Ñ���_\�Tl�b#x������M{�=)���r6���	���Ϝ<#��h�Dm�U�s8�T�����#O~�4��OYI�|�X��˧���gE��̈́��V-�8�gP�|�?	d��o�xjk�E��� ��$��A<B�ӗVl�w����׳�5������ʜ�H�[{���K)~KK��O0J��-q����P����1���
Gÿ��e�,y��ZÇP-Ut�uH��l��=���c�L I��l%�-��
8���u5Y���c-��a���(x�8\	�۪+%���΍M�ԑ�c�\�49 �c�ib�c�+R"��z�
7������šU=-o����S�����OQRg<��-g��4��7�q�,��a6؄]�-�Id��Bt��i��EK#�R@`w�����y��5F���6����|��(�fG眢vF��	kY?�k/~M����+�P`��X|SS-�P�(�"��I�:�<�l]���$ȗ�M,'�VCn?�8o�r��ղ(W_��*W�[�I�w�hi��I���� MDr z	0�E���,l���M~Ⱦ�X�P>��1!��L����>04���JY"UJ>%@�Y�!]fF����p?m��;�L}�h�PL:G����姕[��yW�s̃S�8�_m�
wWt�iD��|�l�mb�Д��=�3��Lʶ,1�k��]n:��%Թ묀:�/&�U�O+P�m�����
AwXS����4�:����
�>N����n�ҟ��OY�F/�������}\o�}�Ȏ��r��	��l�BAk��mm���ڝ@*/Z^ܜ��j
��v����[G��G\�>��->s[��������3��kz�� �, H�a��O,O�'�6?L��S��k�2pө�����k6�����FJ{瑩����X�n�+=��pH)� L@9��|���%�MJ���Z����3�4�x��|x��"�I�j<Ὧ�y�edi��cx� �ؒ&oK��/�!0�&.W�ng��eӘ�0oS�$5���%m�n\�5�=���z��䢺!O�g,�nB`���A��� ��\='�� ��g��-��$���z�D`��{�i	�b��<��>D(�L������wJ�y��6TZQ�%wD��5��g4�/��Y͓��o�:���+;ô��(S�7R�X|#F���(2��ߤ eFE�ه`�	d����@(��Ɂ��1�:�HB��W�� vST �1Ï�klcm���q�8�ZK2b+�)u�����ن�o�
�a^C�����=�֠ <p!^�S��-��LV�ȷSB �ǌ����z �G��r�K�\e�����s���P�s{ˏ`��<Hg� �g�P�}���V�	m�
6��4�M�� _�C��v��u�fE� ܑ���*������$ ��"���r-x�{��� �k'�!���X$RЍ��� E�y�̪��=>���A�n����%�؝#�����<���R��;�N6!�v����I<f:��U�?ri�.j߂��lEѡG�U�# H��O�<��O'A[����G�z?ss��b�y3�4��ժw�Md0#4�߷�����#����\�-@粭>vT�\[��p�o&��y&PA5�R�(�D�	��Q��E{k�Ig��*8Ϝ�r���0x�ZQ�|��@�
���'��n��- nhl9+�C��+�m��(CQ����B���8"<j�ƭX�T����|;Z,�e�M�@�g���#�WbbM��F
�`N2��K��Y�n�:4���.�c�v��DN�j�M����𚉰��a����U�j�U:����/��!�| `m%1�+�(����{�rы*5����/ ���������@,�p*>ѥ�(x�X�5qJy,��e���-��U*z~�b��}C�:�lF�g�Dw� G�$#���7�*�h��F�SQ�G�P��˕2JҐŁr@䨝�eD�U1:4���f�@>��P��$�?�p��wE��C���_I.��pK5��y��G��<&:�OR%�E �Z��C��8��=�_߫d���sؼ�3f���u\A=Ҟ�fX��!���3�=�aص�	��u⤙�J	���AE%�LУ��4�R�:О_h�y_=@��M��:�o��m�}�so5��O��o���晜CC���rha{�tz9%d�����N��Y(u�&
"1ֹ�o�>NhT�Q�t�u�\���e�F��d�v�H�v�w��;z	o:gڃ��5����^a����eTr�]��o Ӌk��l��tГE{O�.��O�L�\�K`���H^�?�%\�^��o�9?-qHp '�Vp�|�(j�5A��a���(s W�7�� a�V���D��	<q���3⎈��~p!u�m�'�A�(��l���wφ�;a%������� K���&�T�Q�6���58�'��0A�-�g��@�X������f9�@¡��K����e�2�(��*��,����׵�� }O��ROjN�O�o˩�'�+�mF�����$�������)�S���)�=}g=�\����\��v �7%�?�>� i|����d��K׵ u'�`��]Y�ѓeQ�D�G��%�G�<��L{�1j8��!&,��D���b���Y���r��fܼ�����ܩQ휇��c	,쯒�9�8�b����sl<�zl9�"�� ��D�e��{W^����,H�]��yz�1h5���m&�،j�7���"��vM�Iq[��XCy���Ö��N[����d�J���l����&���I^O���<�E9Mz,d&AP�ى�O�=�+(��nj��1@�����i'����&��̜`�a�h��Lt�#�^k,N�iUV.��f�D��BNul�w_��!x��<p���b��8��G��N8�#���|�A�s\�`��PW�c����\���ڕ� 5��qP�ݞϡ�R��m��?ZF|��ɒ��
�w�m���1=2_��Y���e�Y$�Z�>3��������Q�&nt��1��F��E�;�ʗ߱�9� �7�3	ԅ��B� \��b1�v-B� �^����g3�!|��M��6P좄��~��(�/E)�9�0@�W���R����9��#��Em����%����߂�6� �W`P���V�2KIx.F�e�0��:7FW�P�T=w��kfݠ$�x���6���9c��+���u��!@$�����sV}�R���׀�y��)�*���V���ю �3B=cͶl	�<��(����_��������1�V׵0�DSw�qf��J�m�p����S��nv\����6%n�DJC�x0=q�u��zZɱ���{�U�#V�����¬o�kTY�X>�?JX�� !�AX�Dd��V�Y�I�C�k*��S�(��ɴ�a x�|���Ua���Zqx)�I7pY�.��<�Y�������f��Ȍ��W���$��f��V�q�b�N��ވ�����J��YM��wU���F�P�#^e3�I�2�
�J3/��x��!���,�5w[s�8	ӂ��D�,�l�Pr��?{�BLl��O��w�'m��L^X,�P�G0�/�}Z��s�����(��0�s���
/�do>�-;bNG�iA�]�>8���[��^�
�F�	����k�"��jN� w�r�� ��}4<+�K�I�n0�_�'~b���EFj�xG�Q���X����U���j��qqZ՞,��Y��0������r�1���z�"1�u4�]�n���tH��_�#g
�"#=-ͥ�;�4�|*��8�Z��%-��t�UC��M�Q���$EZp����Hb�Ll�_�bL�TU���ts����	�q�Wx�|d/�(�g"�!7`��ch���F�`^s��j���;:ƨ��pgrW�T��Ya1��iT���ؼz1���N�*����F��K_��y��8�=Y�~�ebn��'��S#��" fz��%�[)`�%,7��;>����Y���;�97�B�\^eC���d�X��{��%R�h@A�){��;�^�n�
[���	3�z�Λ"2&���"?���ǌj'cDA�Dg���,�Ai�Pk�iPV�m-(��#�s�R��H%�zV��A����a�R�>�Y�Iu��3���N��?'�Y(�?�+��=� [�����v�Th,�og��_j��7��V\�����^���?�YN��'���1c>�?w��,�ߛ�nx@[�I�q�������K�j�Z�$B��02�bc�V���'{>Fř��Eq��.}UN~X�4��F�lu�#)�.����NC�<c���M�0x�'�n����J���.L�uyCh��p�b������1����m���o�9jF� Ƿ�)ȴU
,����L��MoH�
/�U.�y��[�b'�AP�_r����۲�ӖE�MKZ�)i�ޱ�$��X1t��3�D
x�;zg�!Z�.T8�3���3�׻�� ]���E���eӌ�߉[)ԅ�$�%8�r2y�ʍG�6��?�q�4�z^@G-q�H?���C�J�=�����Q0+��|g&jP6�`Qݼ����^ղѼ��ۣUi��  ����B"ꖔ�k��(�`�1�������(lj���%�4�����k;��e��@d1]/���c�V��u��/X���P���i%"@i�1�\G�K���~y��d'���9		����s|��U
GY��;�Y[��.�Pue
��Iv��ѵǋ�_���.��"��;{��	��:�8&Z�r�{R5�p�C�I�VK�(�ѐ�RB�|E����=�_�� �V�ëZCT�z��s�����F��� aÔ+%m�<+�_���8���4;x"x.4 ��b �`.|�T)H$}l#�>ݬ�TOcѕ�������@�:������S}ٗ�bǑ7�aF���N�F��/a�� az ܙ�9̿��lű\�q�x��ad�l3���B��?�c(����DyH\�j�s򼲳��a��Z�ǥ�d7�dBx�����"!��Q*� +9���\�D���dv��DT]9#�b�n39ړ��k�w��c� ~�G<1ǛG�J*�Ա��r�ʝ^����nWe�o��Q��bI6)%�+EUpHb�OG8�%Q�jsꐳ��S�_�yE���gL�5M�%�� !�kÃ
D�$����}�;�,7�W��' w��BX���4*��c�MH��ۢ=p�h4���ф����,��Vx��S����}�b�����T �VŴݎ�i�;��@�z�,��aN������ �P��X0?]��A'e)C����]A�F������L �5�b#L����e��Dn�'�ǌqw������1�S�����bU�B�S�y��2.���i,P@�	�_9�~��N�6��e1
.����y�G6茼f@�<M~I�MI!���u�J�E���~}Ң���:>�ύ4}�*�Ł��k+�BۆӤ�)��<��ݶ�Z����o�n*�����2�X�r�g{��ך�m�(��O���������-MlFԍ�1iGey�q�� Ɍ��UX�Ի�b=��@�!'���Ed A�Y�+t8���7�12�+��8����޸��:Wah���&�Y����Lj0� �q�@�J���.�H 7�9�͇���N3�
��҅*��H)�m�B#�0���0l�J}�,k,��(��.�tbx�]yB�BCeQS�ђ�;n��dֽ<�\'rV7I���?�!'Y.=��Ӣ���������1'_˥�?��j#��KuI拄�J6�%am�s���7�:�k�� 2PӞ�-�0V?���S	�1�)�l�LH�q���)�R$�r�^�H�t��^� �g0���R:�ʐ�S���}�K��J,u����[Y�gK�y�٫G��0@*�-�~䦈�D��>;t�͉aa %?m8��xl /*�0�s�7��r�5o�t� �Q�A|�N��cBL�Vԟ|'�S֞|�c	e$�܀���xY�[�}����.�iC��ּ�������S0NA�J+��4`��:mE���3�-`49��3~|:2�F��N�ы���ǴE;/�?��/��q�]��*{
p�-�,!\��(��%����B�XF�����,�I���}�[|/!��4+X�.�o?�����8ƃ���隸_9䠣���L(:�LE��z5�J!�Q���p�6�!���F��TgΓb����L)��4p:�_��?�O%�(L?�6Ջ��X]ly��iӀ%:F�o�;��<���U�?�5l�E����8'�7�d���ѱ�G�;�}p�<ƚBܟ+jĉ�A�?���Z�\]A-|��<$� ��	fj��b�_��x�_^ޜ�ۉ��d}8��I�����8����v�s�m�aXV?	�i1NE鯫c#�G�c?�u��u��;�$��p����D�ے�xԛ��Rhj��x�ͯe�)62�
�y'��ח����să�1f�!ڦ�T;(b�-�k�>Q$M��i�
����eё���F�m�k[�m��d�I��χW}��09��>�а<u�u�"�k:�eR%����+�XgKw�s���I���Ѧn��Nt��9.�Z��N��ySi���b-#�O�ɺ�Ci�>�}��C�-6�V;Z�f�����F���N�B/�㩟��].�J���<�̠�{�x�����
����U���g �]�h��D%\-p�ٸ�𒕴J5*��܎�sI\�)��u���G�(�a�Oo�P���h�t���q3����
�-h�'�K�ӂ��&W��}�t��������O�����g'�.|��ǻcs�uudqf��BOO_`Ue�Ñ��,&&��f�&�Ҡ.�9$���/!P��:��n&���i�0g�I_�������-�s�6$^�A��k�V��ߧ��?��4��åu�d���P}"�j�>�cn8�W��V�����WfC�QW����hw·�̃��d�(H�_O�+��X�w�1���J�'��bM���,b�$>i/!
Q�EZ�)��v�~s�=�b������e���)%E���{��_�x����r��@E�㼲PQ�=�>A���М��2%3��XB!����SOz���g�&�W��.���T���Dq9�:�|B�6�����I�`�I[[7d��J7�a�i������ �\S���?T�����α�)8ڨyWXAE�D�_j-^wƏ��O 7%�H��<�M��MK�k�I�@-~,�M7�k����*MfϷk�S�bn�Hi�t��wB��}���ɪc[D�+�j/��j���RC<#Zw]<�!y^��&��GՀxgj:8�:K�}|u$�=�``G�N.?��c�;�.�Rd�����F_�:�r1@�{���M����P��=� �p���a�A�y�(���;vP�r2{�q�IG$Y��ݻ�&YTt���:���yR�l������*�[0��o�9�)rځ���T��n�܇�L��ǟd�HL"dY�7+��+�	z���g^v�X!C�=F]N}'z���������?��7�$?�ՔrJ�V�n�9a��eo
vED:�D{�
��L��;mZ����Q�!4�p��t��D��0��R�E��;���	4�n���6ߑ���3�g�b˗"��!s��.���>�.v�c��z%�>N"�$�>�U!��53��������]���$��vƕ=�0o~-�ω�Zo�on��=�t\5��/�"0�#�E��;�����%B�%@]�#IE��!��A�+�z+�L���ި�ݴ�m�ѬR~�2x��#*��[s������-['m~Z�b�����f�#t-����ږ�
���<o��3W�]����1"�����D����,h���.8ٯ�^j5�t.'�p�F��fݽ�����]
�������l�	��8�!;Dm����El����3;:�w��\�c����]�վI,J��a��s�g�L4Ɯ�2�r�y�T������T��q�L>S]!ӧ�0���A��gpt:g�	����t,4k����.�K�yY�C,I�/Q�Z*�b��<�m�
6�π,�x���M�\V���=�;0!���0��%�f�i�H,��N���zP�P�G+"����V>���R�����L�>�l(���9��XN'U}��$�w�j���f���ʘu�^�_�P��qK���~�i�hF13L����;�=��ἷ(y�W�D�nѱ��Y���v�!�j`�#���::�v|I��{V�"h�����M�x;_�ŋ�l�-�O�rm/P��k�v}T��_Q�'����#�V�#��p��6OB!�I�{W'�K�,�Ð�g㣪>p���䦖��I����p�؊{����m�r�;Kv=�ـ
��P�]p�i�s�g���H=�;./���(���i� �������:{=~��&��y�
��x��aZ�a��	�LTtV���E�� �z��h �҃�Jtr`P�̒ �L�U��	��o�i=4�}(���b��D���γT�K�E>���ߙ�	l�#d�+&;�T!d�P��M�zWGe�<��ɔʝ��\�D*R5�J��p�%�3G2�\+��C���x���[b�v<He�ݜ�?-���l�c�7KB~c�f�U�!'�¡r�D9�Q[�*��E��wqd(=hX\�S���9x�y�_� ����]�i0�#S�x#5a8���c��e��@�ZBA)B�U���#B%�q:H�_t��z��o\���,4��u�?T�Ɨ�T�4������Y������ѫ=:�8�h�./��Hƹ��އL .dL$zخ�T��g�y�"�<D9�B$��ۆI��Q�����YJ��u��L�thb��3�am��V���H��n�/S��pΈr���&f4�H(��]n.'iŦm,��=nˀ5�0�ꐾ�H,m�%������1��񱃽���[�$;�|�P4n��%c��U��5�����s�A���AM��t�ޱh��S^�����ۘA_�a�x�ˍS�M��s#�O0�����?
��_���?¹7aa��E[��~��ơ�W���� 9P�����?Y���X2��u)��v:���?�"��|����n�[|8�@	�m���n~V��Nlyi�; Á�g�gȂ�ô(����v��z�]���L��H<������m�/�ɧ���
	�>N���L�� ��)|�W�T7g��N���;Z.��to����;��6��5)�wȎ�9�����R�ryxJ�� �R��w�UF���x!M�R���I�e�q��}lF��jp��C��DE�w@T@6���Q��Ď���G�u��n}o��� �5�'���T�'ʡ�����] �>���H3<w�uP1�}a�4�o4#���O�h���n�A0m{�b ��		����@h�!e�������\�y����T��J�D�;|K+=y�RL>g;�����m@�����?a��=ӖM�JvIB3��sI"G
+.�������:������r�fۥ�ϰ_4�!�O}�O�q��@7��q�V�v��v���v��p��������Z��a�o\��T8�٬j|�S�
���D��x�d����I�����>���ƈi��&�G��x����K�@(�0+X4":�꺞����0�&�i�
r�},@�(�~�A]�D$^���-�)�/�g�׺{�yى	+vu�_����o�ѥaf�����s:�̞��
�����$y� �l-$|F/M���ӐH�0�^,~�Tp��v���!��N�&~���#�Id9k�&�2c������{}���8%��Fn��sy��ļ5��ǜ�کr�5L��ɀ�"J qTPu�6�5��5�8F<6ƙ���IR{��_kѱ�"=�O�����s��žOV�:Ub�#]r�AR�}��1��
Pm�-"���Vtx�q�c:���K
�:Ҙ'⮗^Lb� 싓��i�D�}��?FYޭZ{7�J�A�5^��Ưh�=�l[���ٷp,���~��X�N7� �2[�k�{�-+������Rt8P<0�K�(��\'�m��V�S<[�O1�3����m����ЫN�*Sʙ���>���#�Жnۼ@�"<�QPr���yM���-�e�/�Os�mOo�m�k�A�j[��4�u��Dy�!��M�}��w(�r�d���k��l���JcѤ]u��oݖko}����N�x� #0J��=��S�b�����,dFd	қ,�P�>�Y�6��2ȭq h{��O�j1^:��@h�]xR�#�����g��=�5�3�ǵ�@��sU����'�6��b[>Xe�
���\�XM^�=�*1�r`�9���i��d?�P9����C�Z��9�h�^$�(��G���㟬[���о7'�D���o*���ܨ�r���Z�@�W��,�J+�T��'?ǒ+��J�#�zP��YA"�U"�~��E�l�j}a�QTDh���T�����EȒ�L��_4F�!1�������0`�4iy\n;��+!��Ubz�N�������làHv��G�0�����Ԁ�-(�����fCx�:�<p� )�@���5�J���q�,�1�3�g!Kq�+��#��V��+�$N�ϒ{���%?��F�`{��T�\b��z"��S���/c�J��eτ�L�)@<*u�>'/k�O��K���t��01>�Պ� �YZ3�[fbԪ�v*�V�HV;D��2�����LC��o]�0�!��~Q�)���3���m�)}�C����4���Iv��+��*4^�s�
��ۖ��H3�N
 ���4/^�g7)���o��k/_��e�
hT�P���:��Z������u�N��+���F��ȼe�'!�u�7�F�� �	ν��Q[aHQ�fza�Cs5lߌJ���uX��{����tuY��朠(O�D#�~O/��<�CE{&����~�:L+ KI�JHv���Ps%��Y��b ��U��db��U��+�!2';�D� �B]cJ��d���t;ץ��V,���f�`;�j:��C/��+d$��!��b����*����~�P��X���W�c���З��y���m<�ܶͷ�ê���ֈ�-��]6���d�^�V��,�� ʦ{��{�3����c�8�#p�Z�7| U���O�͗�b���j�/\��B�iRM �	�6����WȂ��41���@�{��B�-&&�b��F�˪h�'�����y%81���n��R�@�q��*���弰��V�*�Y�(�,	~8��״���×�	�9@1�!b9�ĥ�����06�s�Lt��'�:U-�;�:���U���C	��&�����LS�S¼��M{i���~&��AKq�8�g~��=� ��w3���[8R�Y��;�P	��:��ڡ \#g������ �=ׯ��zL
�7;���T��Q51�#�X��V^���ѣy�����^F���*6YBZ q�D��|��^f~��՛��m_�e�YH���G��������#!��Ƀo�Z�M� ���D�'�z�\��Um��զ�Y�7��/d�v�q]���lSU��YCuP��G�S���b�d�y�k1AUk6���(��SD�1�5k)��Z��ۃ��"
Ŗ䏞����x�{o@)���7
�4����h���Smw�r��W�&�����+�jm�C�O�$�斘l:�&�ʏ������-E��{�,K���}�|�r޵�՜�R�U���\wQ2C\4����\�A���R.K)��+s� ����Nrl��"A���W�����ZȣX�~7]��C6�������	� \��H�Q8[�oGx�b���n��e�M�4aOO�����-����o[]��`�6
���5��)���Wd��?��Ҋk2�ܵYK�[��_��@�;Q�szlD��O¯n��<�R8'���Xlp�׽:�Sy�WT<I�E�ˏpn��E����ႇ�#�� 4�AW>�̔� ^�D?���J�����4�����Vk�
>���&��7QHR �C��|7!��K3�*9�� t[7Fon����b��CV��/f%Y׀�� Ő�ªw�w��<������fb�Zx><�KL��2]�B�|�Nu$�F��LRT>L{^<�"�?A��r1�a����`���֪`�=���P\���Ïh���s���*�A�VX.ќ��-ق�LkP���Z��Κ=hyz��Aʢ��/����5X{��a���T�8�����$��@w����tS��zI��ۼ�w�PVM[{��C�8.4q��!.�SAtAZ�jc�b�j���������|@��]��}	��O�2����-�f�`��!�Xg4�������M�w�T|�v���M�EeYz�:7#�z5�U�=�$�����Z�W���#^y^#�� wcƬ�l#��ST:�)�c�&��������ɣX�Si5�
���.`40�����Oy4�P=&-��h��جrH�e�e-�Y�f�|��F�ʺ��1��|��|o �ġ6i��x�;���֍ �� ���HU�WM���C��P{]��@8	��N�a�aU Kc�h�5��Wl�}����,�j���)��r9	!��c�Rv'�[_�x�,�kX���r�1�?Bf����1���N�À���P�քJ�B\�o�ԉg޹oc�Vz��� �j���C'�����e�ݛ�TD�S��
��@3�����u����;:G���Taң@1ʘ|ݷ/[�Ѕ|F0���c�
�	��l���n�~Dԉ9KgA�"�OHu�n%oW�*$���騚�J��'K���CFvUi����δ�kp���9�W6uǏ�x��2ػ
�?��.����S�mn�SJ� �ܞzο�8ʇ
n�~�cͪ,�7�C����]�.J�l0vjBT�A�� �j�/��L���/�۳�J׭;�n�L��T�i��ft$B�ͅ� ��3�v�"*��f������A��X�@ +�08|�~��s!�Z���#˻������,��;���E��?�e��[C!m�:ݎ��!7�l�!��1=�����\z������.�� �����A�%�ے�8�-z&W'����k�ծU