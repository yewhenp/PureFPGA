��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ���\::����4v/����1/�C�s�d�ǻ�Pf,+V�`sBo3�����+��AE�YeTUxR{�l7�eZ0}{�믘�Y�f��k���X	4)I�s)�^6F��?&�����`�l��y��<����h�b���^J���l��2X�+�Y�IuMB}4���.�~��a`ÐH��̳�y��A����05���ޠR�n�
�OS�7��FU�J�!#�VZ
ĳϴ��G_+!��h��-��~GmGi�T�g��
���`;(��/'%�>U��F�g��Xmb�Aސ�;}�2Us����0��c��Uk+�GG�4��@8�iJY��Q,���.t��˪ס�jﲡ���e�%]�V�ٜ�x4sa{����ܠR�vh1=M���д#7���+�ϳ��N��N�	TqU3�n)�>	c�\c-꩎Lu��8��igOk����А�;>7j�ط�ק�!W�7�[�e%�G����b8�.P�A8�yr\z_�OC����k�vf����/[��ж�6��o�j���W�0���
�G��#_����2��d��0*��\6"�JBv�
5j	ؔ�y���[�=��_]�z_�ω0|~O��2g�~{��B�f$n}��hI��k{ au �'%�ӏ�t�ѻh�Po�vi�
ʘ)���s���,�E��0��+'.C+k�\/z�3$�6nM���p����커��DLr.�)<U��y�-X�@w�u֘S�#�n7
ѭm
�������=_�Ш�CX#���e����dE��D�ý\[&m��o�\�FSXZ��[`�>��\-IgQ�xh-w����q�R" J��h,��b�O� ז4��.N�*�_^� �[D��ŭE!ʌ�ނ+:׮W��S�����:v�<�׶��}�p
2[�j�k_��b�Ϫ`�MPI,w�]�^Q�l��(o�ø>a#�~�ɓ?���iso�ۆc��6DM$�"��k���� &�n1�prӾ�rM���Bp4e�xg��-����1��RA��F��_��m�?ڥ��{���P�-���nH��v��>���>IFP���TX�~m3���ԑIz�J���5��>�2fm�(�֫J�� ����.}�H��<^~��Z�����QD��Y�i�!ʽ�./��Vd� ����	Da� ��0G6;�2�nV�s���qۘ���T"�0�:��o6�P��_E�T" �xT#q�~
+�a ���'�4�X�sf<�d��Ȫ\g5��?�� ��4�O�-b$�1����!~�ץ'��~�Iu3i�7'k0f]���;��V�et�DkR�?4�I���LJ����K4��I�F�%
<��~�� b���|���W����~ECm^T��{�cjz=�J!p�od�K�����N�� �#��@������yKD�C�K�&ItqH3�P���G�Ӎ]��@#[��|��v���Z�@`���b��I��RƘ�:�
9���܄g�g��͟�v#9j�9�ً�S�(�}���f'd<�Ӕ	K�!*��6$�'7|QWg`mX!g�B���qGDYk����S:?������	>f"�H����Ȼ�������w�k�������T>x�b�&O�r����FB�w��oC~��]������xg�9��b�X��z���=5��8���u�{�Og4�9���<G�_0^��U��qX,xO�`� m��xp�;O��s�I���ҙ��%dCO�$8u	U,���m:r��$�o���g���\ϳ������j�U�¤eT���2�?�^���Γ�Nzp�i�~�[�����.S5+
�a;
E0�e_�F�n8����ǩ�B����=xyْ�ݨ�a��ͽ�ȉ�bc�峍��L��b/S/��'������{ɭP��+L�^�'�D�.ݤq�b�'�+�n��a��S�F;�2��%p�@�KE�����y���4R�����{���Y�E��2���	��0p
1w3��R�&�[���'��ilK'� ��\���߆pQ|9�9�Lga�Q�܄$��r��Φ0�pq��T��Y�yw^)`wk��,�u&o0�{M��Ʉ�R�5~{��$1�sʳ��mZ ��%���bc*�F����`8`�{ˠ;=�46�ɗRy�'���?��9eM���I�EY֞�>��?�"�܄%a�i���(�<�Jk�Yݱ�K�\&0�l6���A{��n3!�1a�9� ����m�Ĕ���/Aś���ٷ�L ϙ�;��g���o��E�qJ8o���.v3���� ��O3|Ӷ	������+�&By>�Bd���>���3{+T���OՖ;�M��B�j<r�QI��=��0tf3�VިC��
��u����6�	���q��g��*ˤa>�ث�8�a�#
��'3���&>��)S4kD���ȹ�?������
�1��=d��2�~	�SId�e��)������E������4Q��P��/KBDHZC ���u�����ԋ���
"�W�t��.� �L�kyb{2<+v[�\�N��Y� �?Í���;�.�%n&ʼ��q�zH�]����~k�1ň�4�LD���C]�d^$)=W�}�4|������T��j�5�1��:є�f�T&���7w4���Q�{r�����5S���Ҋ~�ig�	�>�ގK1v�!#	4M»�2sZ�)�e��z$�����~��u�t�}�����Lj�6}��x[�V�2�FB�{bX��K���!�PE��K��� �"T�BM
+���A���v���nu<Kx��@�4H u@u��!yf�׎�c�a�rg��Lu�S������:���]�G�7��l�Λ���D{�X���h9��]��S% ^�A����2�M�H�)H����_P�~��.�����XS�]��	Օ�wS�YWތ,�-s�cɃ���E[���-/O�����G��I ��
��SD���P���Dh�4-�F��ĳ�r��ol�|�A&eM�?��Bvj�~�!=L�'x���q�����c2?�dkJo����y�Mձ�ۤlf�M������o�d��s#�F���y���-�~���
9��ڰ_��@��=�f6� fY�kk�B��k� ���]���Ȩ���{ �|vG�kd��_��f�'zm�+Y��9&�E�2��8Xo��!�ÿ��ةs·�NЄv���s��FK��%q+M�m��q��W�ζ�Ѝ��\�%�*��h�倱X��Y�v�����<m$Z\��st[Ƀ��
�ZXB^�W=�ʣ�x޸�������= ?FM����a_�vH�<�h���K���G�L��v����c��;��O�2͠�d�9�.Ps_�F�ӇfJ2�w���.��(�:d�d0_H�i"X�5������I�⯬ao�Y�>�l�[q��F�V ��IP	xZg�:l$��5NOۛ�4�>�A�QT�3��5T�cG���ps���!�Ӆ�G��J���K,V>����c�7�A+�BG#ap�H��
�j�s'ԧʈ������f���$/uܲB���$��.����7����b�_֑���<����B�і���(���AmΦ�YX��׶ĺ�^6�qգ�t���!";2�w�Q\�u���Q-�3�~���^Wi�4�-Kۓ��! #G��Q�=6M�d���*�Q^���億DY�z�&�}�U{��G@�!|��[�
���7k��p��h7�&��<��`Lk��r��Q�-�>hO�*�3�*��b�A�6B�WY���
�%,7���E~�5�8�e��K���[�yE�Y�L��X��tTE�}5P �L�3y2^X����\<�ř�,+\��e �Cry땑B�T5��,P�U���he�s%�nTw?ú�	&�:*yiNA�Ni2�g> @�e��I7����.t�=�"���#ǧ?�
;�)T�jVз|?�Z|)E��#L��$t[���`Lؔ��P��u5-#X��⏑�९M~�Hy1�6���f�Z��i��_2����mW�ĺ\ޏs�˟X��ȃw��uz�[�F���-$ �p�j|�;6��x�v�Q�k.�<s��TDT]��Er��I��JVX��=����np�M�b��,�.�v��~��p���h��&�-����:� ����k(+ӝMZЎLD��2�{I����ۿ��+�+o�H)�gL���'U�2-b�U�\�ΞΈ�Ǉ+do�4�ꈀ�
=�&�B��G�2G���K���fb�o�wA���_ap,���8�;@�<ͅ�A�P
a^)��c��-�vcjr��fv��T�[3w|���eb�~H�2�y�1G��AG��3�}��瘡D<��\GVZ�����n�� :�T�.Ї�'��C�y�̢�I"}��܏�*�?����P~2�U�ϷyL��ǹ��[֍ھ����P���p��Lu��F\�S ;4Q����6O���Q�N
��1����+�{�6~�Pkꐠh��eL�Xu#b6
����%��6�+NN���@^�e���[A���S����J�8.�>�{6���J,{������k�o�3"B
sM��:o	� Չ�E{��*؁f���{�G.1T���i���8v`!w�*��Mk�k8H�E���Exn�1@ƪl�K���cLx��*�G��r_$�Z��+�{��v��nyB�
!�F���%uXw�h#6�u�.���H�dquq0��l��>W�R}�s/�$�~e%Ғ�i����p��\�HJ�_�����Ʈ,�����R��9v�Ձ��w�ע%��k����3���%2���lw��������|�v��N����
��(6;<?p�!�!�,��U�Ȭ���Xs����r���Z��0i�p�n0��V{��9-g8�O�,��zs�#Zƺx�zPYZ���h:
&��f��c����k�q��>�4��,�ټ�����a'>�)ڔ��ԩ_�-ŝC��c��ɛ��r���
��`�A�*pN�Y������;ZL4a�0�=��T��'���9sֹp�`�b�lqvr_Nb�cY�·�4�S.�X������'�;f�;��Bg�ih`�>�U���a�r��=m1�ۚ3Éy}3��(�hJN0g��֜�����^C����i�t��h���X$�ű`CM��H���,|�yGh�@�Vco�bNh71��G�T���Tz�F��b�[h��v!�m�[���B��>+nTN�}�GZ2d��.1K�e�`�n��ǰ)�H^ܸ�_��ͺv���ª��~L$�+�1�=� �r���K���}��~l �c$z�����"<�*��N�m��7��u�7�U}�u��)�����&� ����%�}��¯�[f���T��/�e��E���%3��n}�r�I��]t��Q�H�rt�9�/�H����SsfFQ��U+�'KtFEq�w$E�'�� ��Ii����v���u�	ə���u.��έ���'���������zC��Ԡ8��3I�j{���~��z��y"�B8$�H�]_�#5ZY;�y%*}˜YëJ΁w�7�2@��$���^��)��P�XE�vEbu��s����>�7"%����ۙӗ��h^L�58P������o�\���=s�� R�膠kH�r��<������pbċ�Ę�0>F&�Z���3�5��]���0�qȪ���[����2� ��QO�Q�u��IW��{����n��J!;^8��Q��Kk��
R�����1�}O��j,�_���Բ�d
X��\���h����Q+�QQ�a��jD�>IB}\-����L��������|��t��u�є�]I:)��5r4�|�7&���ƮcPHJ�4�]���Y�8ҧ�_�(G�R�^��$�6�s7�k}߸�W��2 e����N���*�`���]�=���6���A��"櫶k������ �Y6fa��7߅pg�б��_�����r��U� )ߪ	E�*���V)F)t}vAQ��1Ɔ��%K��{rR[���œ��R�������x�*��gA	ɇ�h�F�&I'
�'�1;��ظSk筼�+���W�ݼvNSw�M�F@+6H4L�n������{��|�i���7)�x��P)�<�����`1?��ԛ�B�h{�W"��Eٷ�A�M� �2C3�AX!O%�!j_Yny����(ڞ���I��%I����l.�+!e^���5���W�1}��<���t�q�BJMڑ��ܲ#��{�xqW�=����hh� I%�[��x�Z -��|t7ٞ;q�%)赻�hdo?NX��ݨ@��h��P�Jd���E��d����PN��Ɨ�r� 2Q;�'u������П���+�"I�\J��5�_��E�k(���h�xx��B��и�nK)[
#�?C�!����<�c�O��Q%�ǁ�B��Jl�� Rм'>�9��L������+(�@���m�(UX�r#��ȑ��n��w�ҷ����J�0L�	�z���pW��P��R1_����!#OEV��3_�O��M�1�STm��v�~���wA��ӡ꒲-D=�|>Ʉ3�w�U�O��D��ۭ&o#Ƃ~�k5�+G��#�q����1��?48��<�(e�58I=����Wcy����2'��Bwy�h0���n���� �g�JO��p���='�a��T.����CHg ��,����W#Q���������������{3=���K�����p�a$ъ<����,:��O��+�)�Z|�5���Iv�%���^Y1ؚB]�]i{r	��LG���|(�/�}	�V�)�v~����\��Yi�)>�F�Q��0�����A�\e#�G(�_g�_����G��$�RU�9�H]�k�Rb�6�ʯZ4)���f��:��
�$�h�t�V^�)�3�Z�71Xb�py��l�g�o� ��4-�SU�1����?:��´r����7��
F|�Qq�f�#4!Tu;���)�y8`��D�u}ާ҈����_>�R9�l��7��!*U��M�et�p�-/�b��	�%�)M׈*#n�A��)���p`h;�������?SD�0�E$�7(�ى1(W��̲�`��.�F���_)̯��I�M�S=�PfI6kJ�̹M��) ���.��`�K�M7���H��/�����QT���=a}�sK�����B >�`�������e
�F��	6��T��#4��LB#jb���U#��q��DMU�w�q݇ߨ�A���x��Ïep!�c�)� ��Z��!���<�L���Mr+��ݲ�r��	Dd��t�f�b��d�!�7� .o�ځ)9��j�%��¸5�9�A:W�ȐS�����ZgOT��Q��-�%ɾ$�oR��Jy�3�-��`jU�[�Hv/�?���8rh�����oz��t$ ���h)�c��v�qIʳ|�~�Tu���ʸs��"�tm)��;uMp�-��.�W'�|��ABp^�Z|e@�y�S�7���A���.ͪ����"���ޒ�;#7ZΩ�g56v�%},m]��P8�JO�W���IP��k?�D��85�B=���0"�1W�X�ө�g%*�^�#���M���c�r�hi��;�W�l��vH��Jfk��!b�S��E�׌ݏ5\�"�"�s8��˱�z}B�0��u��L]��`��B��Ī=�����"�s�I?�~H�c��3(�8Q�m�[��3���	3��[� Gq��e�T��/�)�\Z�,q���8md����S��:��~+��x:^�-P�B�!+"�'C���/%c5��-!�s�z8a�����{1���Vx}�7�T~�=YQ�9^M;R
"��Rp$�t�$ɴ1�Aaq[ $�	�H�b����-��KJ4.+?�J���U˻��'�x������w�	~�)�H���;�t͑"�-����p��-%��c�N�!H[�
��W��CGٺ.�{��À~�j�oA�Ë��s5�I�N�7���XXU�@�^���'�m�\�:�i��پ�J���W�,9Ts��u�H��M7���!@�&�,���\�k?:'�߫,%�,���q��@�?|'d�tG�i�>7�� 4��ƪ���L��s�<:H�U���»�nΗ}�h-cI2 ��>%K��G)�`콕�Ց�l�M��1��HH��Md4�*��D�W�Uc��5p�{ў�g"O*{�9� $6�H�zM����Y�GyYAT��=�1
轖���p�gŨ�S��1H�M��h����qOwl�P&/y�\m�tl��W��aU	�/V�g
^��!��A���sBA�,fw��h}��V!X��n��8ԠdXA�˻v)J��{ȝ�Cz:��n���6�	��n�ٍ^^}fmF&c�&�v�Љ�+џ_�q�[�Q�]U�g?M�̑�Y�����]igRpLt6>��%&�^��@~����Jh�~Y>\=�p����K�-�T�$�Lpc@�P9���´I�~RS�Ŧ�����?�W�ޭf�%�M�D�h��K��b@3q��I+04��-k�m�84**���3�"zoֶ�)�,�g�N��v-�p$���lf6"��d����1�$�K�����d�I:Pos�P�S�O$�����#{�lm�}Ś�~�_�wF��a������£�{��CN�Ղ�]�.���qH�(�==
[���+��Y��)���Qe~�GJЕ��Bf~�|.��4ڧ�)tϟ3h�8���|\S��$�+��`�C3�>��k����O�f6̎��yqp����}����OC�U�������ɓ@�Ί],�ɏ���(&��Y7���~G��]HSĪ���?�����?ȃ�C�R$�D�/��Bt�ܯu���8���V&�
b֚��OG}��sG��>��=�5��R��%�wVO%{�6���Bƛq��-jC�5�_pr ����U�;��&�L���zϥ՛\���#�T"̿&6ܕ�8޾�jk�Kѷ[M�)E����'������<a8��[� <,N�n<Z��N��@�x�As��*�����sU,���0�Ha���\
T�'%�/ �=�gܝ�0+�dA��x��.<��	��&��:ym#?C�Y�7lS���?.������U1��%����1���$'N����y�u�.G"�oG�m�2F��:<mH���k!��i��BR>�n�^5�}�w�S�l���\����b=�S�ae�}���l��6H��ER�[����1���B�Z��q�w*��[:�X�׎Bk��Hz��蝬�l�>�ٜ"k	?���	��<��C
Z��W\�:p17���0���'O�50O��i��[U�"�E��/�qf�<4gr{�k�����i	g�tcY����\�{Z�����kছ!���&�.�7���}��*f"GقeN�	���ܯKD�T�'�T�ȸ�~�����s���E{�M������G8@Z[��7]���)Tp*�zkk���M���0�%��#b�U���:^��׭��$�"�YL�;���j�M�7U��h�͆�0��+7_�V���nq�=�����	���x� ���o��A�}� ��P{׈E)�kT����ؗ����VEw/��Z6L8�4�)Ǟ�Eiw�F�wW���;RJ�a��|�.�G���$�~S�8/#o���Ʈ�.8��UOaQ͞��4�~����;4F�6<r��G�t�㮶 �*�M�K����M0�X��h�[婗�<��(����)Ȁ�|G�Ef�
�Z��{��Ȫ�(��G9;?����qݩo��ȃ��K�a��NðUy�i��;�d�5u�-9o�۬o%o�}���-Z�u���r����)�3E���_.>�rf���}�/,'SK#(y�q�^��2'��ފ���7��~�#����C�������T��A��p�{R=W$�L�YRfkV��0S�����u8ޜ�z��6�:z.h�Cghip!?v����*��W9�`p�(�������Έ9�u1�dT�4���oY�?2�1�ŹɌn8�JJ�_Y���#Z�۞���ms`Yed4�B&-���r�e���ޱ5=ǭ�Q�}���HH^<):8�G���a
��9l�d͒r;�3!�|�R�f/8	0�N�o�a��>�Y��rvVɆc�� ��!��$�06Q�{���8=�~�l�]b���2)���\E�%���-2��ǻtY��:��$�uP�t(9��v|���d���6P�2~�U�e���ȳ#۝�b%#*�1
]�ͷ�?�Wg<�����������Θ�+��,��BXC)�`�-C�7�.�<(W�
�Z���vZ@~Jb��[���"u4��Ǟ�4��NZ'����	����?R"m�B��ct���@򦦃����:�U)�}���g����W�ꂗZ�Q/2���,�@0�\eSA=#���{��稇�����#��"3b����6�)��f��-J��c�9�t�0�Na�J�����)���ʄ��t�ٱ�����ݝgH[��r	c��S
#�uiU��ei��+�����]��[(�S��vJtr�w;x�ӴZ��a�@d�_��}��?��*��r�����Py�C<��)0��:�L��P�l~���q�XY�P��@�#84���~����wWY���Y��|R���\�8(w��
bp�R"B��1�}�k��G�P���+��C�,l�OhIx���6TNhA����9�&�w�b���'
���Wh��g��i��7�]$B�z�)Pz�/_^�P֪5_�_�|�ғ���H��V.���v�B)ʖ����Z�<��Q��:��b?Tռ�)U�=�]�z/����@Z�l�?`�}T�$�
+L�kp��%,�Bb�d����D%N�s�����F��<�7	ձ���7�w+j5���@�7<!�L�騜ӁVW�cZm��V)t[7K:Ȩe��M�������э�gj�l������Y��I�,�t�[��I�/�N�;��,�4N����ͣ�~�|�7�Z��㺐|G������K���[뚷�g׽3ꂫ
�2L0h�4��� xb�����2Zh�a�4N4���e���b���6(E����he�>P�~\����{�N���c��B&ʾ^��Rg���[�y���Q���̣&A���*�F�Z����zk�C�'=�r�_������3I o-Z��f6CQ}����K\�-|��yU:Z�M����_z���1�&X$D�;q�VMA���|Aċ�0V��+�y����]+�����ϝ+�H��q0HPn�~4"ׄ���e�uR�\ޚ����X3�\�Q�#���e2� vk����bֲ�)�SL���r(J\A��9q{���3�m�
�(�}(r���w��P�%D�\ӆ`���H��~��`&Mk�ę�|�F�C.-��G��4�=t Z�_�/_ދ1�.=@������6�nH����xu��ܣ���W�;s�7G�U)���p�2�ǯ�h�G�����-����5�`Ըw�p���	eS9Χ�u��I��>��k8����+~H9C��۷��j☗�w99��07ᧈX@����2m�%�	J�uT%��ը�Ӌ����~���b�K߱0���|����(��.l!c��4�����f׈�y��b<x1�H�&�f/��x_&!��S��O5Х���z�e+Ҟ^�rE�&�3���v�j�_��<(���G٦��c�O�&b1/a"Pu4�F�cզ!���q(��/'�S�n����>���xP����l 8A���j��d �CKn���Q�]7eV�Ym6��i!��/3li�g�>sb�Ă�=�s�8�|-\!�	&�ʟa��:�=�������I��m���n	�	����iF���M��D ���mY�~&��e��4��@���=w���۱�x����8��x�q�^S�`��[&v-@�rV9��Z�kr����=���p���ޅ���#t�O&��O����n�v%q��V� l��&���X}a�c�t���
���o����X��ZKÇw#"�.��㹗[�H_c~�O���/JuH���~����3�9�fR*	>�ǁU73x+U���ɑ.��&7I�cri!(���@L�@�����XL=J����W)�l��n)��3�/\����pR4.��Pa_�B#�Ʋ���H��N����+��`�ny�)�+���{ې�,�2�0y�W�?�LrIӨ��6�����H�=v����t �ǎ\��^WZ�^�����W���jm��}��u��Q��,�d�U�{���f�s���ŋc#̹�S�ȓ�j����N�"��42���R�芚Hil�`���D(~}��E��?�c���Xl0���w��>D�cˢ�z*S+���u��K88��k�hsw�n�&��;!�1�?�!`�/$Ic�Fl�ڸ�;|2&�0k+W}CI�e�@[ҙ�������
p���T������x)P�����X��
�@<M��uH}��)_�-� �W[���&����A��]�o�Iި`��/�\Ʀ�|x��|�N �ߕ�_Qz��O��f���1�z������7Ȣ�Q%�m�!}c�J��m���0�}\�xӴ!�j��H ���l�|Z.��r��>o;��"�GZE�0�B�a�/W.�-�[�y��]���O����G���5s��5��^�aPg���.�e!Ϯ��JeW�G��;���$��yv:ۦ��I��C�(H%��@��,Q�������	 Ȕ�
�;TRS�V��\�+B��٘�':�� V�s_�"X��x|�K��A�.��t:cLR���(�_5�0�����1���x��>4)@�m��Hth�DK����6��0���'=�HB0�r��/9�����O�Nժ�������5���_vtw�0�F0tJ:��(��2ОG<��nc��b��ғm�D�b�W�����0�.&�E��Y�(��h7�/M���8��ti��J��k:z#��2�]���ҁ�$��11*�L|�+�MYl���L�����2��R(w�ue1^�3S	���9�0}�������-�g2^�R��4����������,��j���Y�C�WH-.>�#m��rp/���� xprU�L�7y�X�S���H�V}Cӆ�����oˤ�\R��aQ�.��L|S��MC��n	e��y6��%�7�|ʜ�� ��ꅮjF�f��J7-c��٧�YC��Bu��X���ʮn��❮��2�&z���o������� RD�5@�I!h��GY��jzw/�6켮;�pC��ʛ��:a&}Ҳuf�:#��o_�[�i��$�~H�g�xg�!����5A��
�س ���_�$
'G���?�4��E����:�K�rKXG"�8{��u�tp}z���X}��o-��,�f`6�9ƟV"x�P��҈Qd�ZܦQ��d�'�+�5��3�b��mvq�=�|��'�T��l��|��'/���9�P���n����f�P�"��=��F����r�[Gn�P��HeX�_���@v�c�������i�) Xx��&@��q�o�S����.Ǉ��w}�����*=v�_�Xg��2�%�4�<EԐo�u!3�D�rU3����3��feֱ 3�,����PA	�sU0��;?�#g���cs�����[2i��QM]�������m��]�R
�=�+��{8F-j�M��I!K$ۊ(A6��� !{��;��0�B�U� x��k�bl����'�;O�0�W��/��S�Z]���[����Q���!���_epG����
#8�/Ƽ'O����ϦV$����/c]���O��.���) �B��A҈�9���,����P�R�P���I�H�	w�1����f��,>��}�N$"ϵg6�BZ�9�<��wz�a�F]���W�$:��e$j�v�9$	�B���L�~�  � �>�2�[*O��s�ʊGҼ�C���T���ԟw젘�Հ���t��_�O����z! a�م����ݎ��KX��z�z�Ó4���:�E�_�Y��&H˱ߛZ}/��[_�b�`r5-��"�pȝ� kS�j�ԃ��<k<� ����/�V0�;��B�O�L�XSR��@���U0�n�V�w��׫3�C�A~T�ƃt0���,ϋ��~sf��k{m���(���pLj�����q�H1�{g���Y `��T�h�֧^�))��BCC"�JB@k��B���X)Ɍ
W_�������V��Y4�.��G�5:(�2��2}�N��%>upm���̴�J/ �h0qp
\��/�
A*���"����<7$h�Yo6i����Mt�j�L5�o�O�q�N���/)�p,=h!�DH��jfKt���=?��p1R�'<Y�bHB�CIvcz�4���P�v�X>O�q�9��X�� �(2�U��0�g�T�٧��^��t�!G{�X@�(8)P�k��D�FcƾvM�'Wg8���W�7�3)J^5󭗬Unj�*�A_�Y�9D5
;��C����f�JJ�JY��"[�rv�ҿ����w%���N��N�����y�5���f��KiT	���S�9��2�݊���V���F��t��'_����ѭ;��ݪ5�`�$�$�@�CX{e�����Q��
�ʞH�c�0-�;��L<|�bW���׬�(��z���w�����3�c��}� �S��U[��?��z��O$�%�@�8B:"7��Sv�	������q�D��Z�`����+p�_��V�d�DAHͱ��H_�oZ�Im�Oݬ�g&D��KI�Sڏ"��N{m�>��Q2�q�1�*�>�B\ii9���vĒ<�8�`瓾��kg>&�z��QX��A���_��Ey\Qm:��lU.V���e _�݅Ϲ���n֗��� �A����h�nd�]c�ľS�!V�w��G�!�
��C!gZ?hM�{x�f1��-̇ �>�K��2�ڎ5���";e�˝�Hz.(޿��f�o���()�Ë�q���������n�S�٦��?���O:}cr��Z8�䪜�l{��H&Ge0�fG������Xő�}�R+��ɸD �Kr�����O�qi�6��`����ܬ_!V�/�J��y�O�����J�t��+�B�����5��ʢ�R/N>g���85:+�t#�s��2�r2���͟����77�7��;���z-�r��<�.��ݱN��S�1��S"�s"�����fM�R�m�?�V�n���a�?`zs�m�D�n��Ǧ��MĊ]���������ǌ��D7�何ջn���ި���
��c�u:������НD !(��^˪O���%�"�\������ɮM���{��V׏'�<d��]�3}��s��΃I�Q i9�2�<��
�<L<h8�Yz���ɭb%�vB���*��zb7;�FB&ב�D1��(G�{p�پ������z��3fحQَ-����(����q/���=���u=t�= TDq)��f/ӌm��/��5b��n��'r,k��h�_��B�Y��Ԅ�Ǣ5?�w�����b+
Þ>���W����viiޮ�����e��@ ��Z�u�轎�\h�#u�wvLY��H>�u�
�W�'-�Ї4G�!�l����Q3:��YZ6Fk���,F��e?`�9���DJ�K����B@,��v�\<���Y޴y���2,��bF�ڗ���R��\���1D���Y�|��Aa�22��@N�Up͆�[Ɖ o+��,m�C�f��,�^�CD=� ~ ��A�d|���o�
.�|�A*L-Q�ή_��������LB>Lَ����w��We�G��Lަ��<��;�g rs�<�e�#}e!�#�,%�tט���qpWم.|wuJՇG/��H^՝�O<m�q�\�m�� 3�D���H3r�+��Ð7�45�A�ƐS,�y���vz���f�0Q�ͨ�a�J���ho%ϺȾ����0_���i�:Z�{~���O�%�k:���d6(����<qGۮ�H&��� �[�K�R��{`V�>O��C�X������Cc9G�.��8G!�H�̞$L����-�)ơ|����˧�����~V����e�zF�L�%
s�Gg)�fWme��y��bX�o�5���?慉-��7�l��#4C?p6v�h�D���x��̆j���L����Oi�үBsDV��D���}km�V��/f�� �ƶ(��ܗ�̋L=b͡�����v���n��SO0������y�뒩���s��
�~��LNP��f%ʞ��,��[\	���ƋaT�C�Ѵy�Sw^��)R�w��ѻ�>��ipl�0|����p��̐�O�ͶW3�i���|�ڏO*����.BtP��E�,�X)�`F��c���G�<&g&�5��'&��mt�}��Mȕǟ�Bm��;��g���vhi��Ʋg,&!����p�n s� ;�Q�̱��#��(~���ע��h6┇R%����fI^2xaР��*���Y���ߋ���W����9i���"�Ǡ:mTL5P6/J�9�o/
�ӫ;*�~F��r/S-��y4H!C�]9>���3��Μ���<�rR��D���]r'r����p�z�]
��fm�*��3[�(�A�Y�O����0�W��岷�����v����N�i�#�QF9�(���d����{�83�TT���Z�D.o�%���H��V�(�%���9��8(��Tf�$%��1z�DmP�Qtw���?q����F�� Ԩk�g����Wt��b�"��d���[S��s�J$	w��F@-5Ӑ���g�6i��˃��"0��B9�<8�˻QWrs5��˭noʹݟ� S|tb�����+6�8Cf�&ge2Bᰗ�ia�(�$-!D�"~�L׀h�2��';��P!�jr'�1otr�\�-c~ZK��(����>U���/~����X_R}*�����#EY�,��f�˴���Q|[���p�i_`��n����hӠ�c��/򵅝M���H�$��yٽ3EU��R�	�:|�	ϡ�f�l��P����E|���NeSvx�LGj��]�����	�
�C�^�<h���� �)4��ۣU1{y�Ȣ-�i�c��V4��f=�}��BS���o"�ks�>*�#�VH�+ùxn�Z{ z��-z��Ր�)�{_�4#D�O���Zמ0�fnk�S��~���z ZP>���Q�g��`�C��S�%H�"s�ȵR��١���i'�{4�ƥ�:nWZ�O2��4��B\�+Z��A�I�-Mȷ-9� �/U`���&��]3���Z���z���J�s���?Q	�Tv3�\�$�`H=G���!��-Wk2����#b���^�h`E��T�wLla�|q�'Ⓔ�Wɚ+8��-�5_U �A��B;uV?�j�	l�\K[�c�9�+5P���CDg��P��;vtɬD�|��`�g�I�_.�k��Ξ���T��Y��,��I�Y�5t��HlP��d�~��%����r�/@U$�����O�FwTHq"�r|	N
��wڈ��W/BYєL��Q`u��J�o�I])�R��8�j�l6VD�D��5�(�t��t��#6*_ӏ}�?m����f�	\�/����u��.�C;'��9��8BO?����T���3�T����e�Ӎ�iq�_z�m�`�.x�Vjd�(F��!��yNb�$`3���P�pr��_����X�\�,�������Wg$�7vH������d椩_�:n鳍�C�$Gknl�^�)ތ,X�RL�ԗ4F|b�|�^�^�?|d��R>u<s�1��6���?�v�c�M,n�eO�����Х���au�@���T���}"��(@��݁�P��g*W�ʹ\mі����޺�R�Nq6���E�E�~m�y�<;��h�WI�/Z/R��A�z`��@���
�P@�aN27�^.�!2���b���J�q�:_�[Zk��U����s=Z ���s>;ae)�����Rl��,}Uh.;Η6Y7�U�{ ��Wmp[|ïbkdtBd82�;�!w�2&3�O|x
��?�OT��,�/�
BO�b��q5��d9K��_���ҩ�#12b�*�ecPƾ��.���ZXswu�"&�sWL��E���E���$�����\�^>�K)F
(���3�bu@m��"6FJB�@=�l��zj�,�(�*�~1�v��	������:gp�Cյ�rN�X�S�� �a�'��1���~��kaۊkP:��V���H���Wqf�0�`��K�^��`����͕ptQ�q�aA{����1�,�Gt�|�I�M o�F����*1؊eF8��"V��ǲޕ�b��������I��3ױ>���t� ���$,��P�W�(�������k+^'�����a��74��q;�^H.&Zۿ"����p�:� f��3ٴ��s�_d���ݓq������^�����J.��f[�#�K�u;�;wlb	j���Eek��̨��W<�&@O����b^9O�R���(��dH�����>�/nr�w�p�F;%����OӗS��%M(��z��M�u+9߬[s�ߎ�%O�%��&�?�������ґ9��:R�L%���y��o퓨/�\�pb��<��nA��t�)8%��=C�6�y��:��0H-b´}�Y2�5���i���3
� ��Pb���������ڢ]�8hA�T��dT���&e���{N�<�Ե���h��쨞�kA������0��Iv�;}��^�cOS���v�׬�L�$�1L
|M�����:�[/�B�m��		`Dp2�Q���2e*���w��_�+3���9lbF��
;���Z
\��!�;�Q���!3���).����<�� ��[�	��p�b�Hk�/�:����` r=�ƪQ�@�ÒX�q����炰*��YY� ���t�o��Oy��#h�+���^̒ϓ��=�:g�2�KVȒ{��2}�	�a�R	V�-t�=�dkԍ\C����nZzԼ��R�tnlSZ��,el5�:VD�E�q����*bU�;ftߦ�7����f;�=9S�dv�I˦+�Kj�OAw�Pt�n(�8�����t��Y�㆏���A2Y)�]�7��,Q��Ge)?�q�kU>G[��S�P���3Zbw6脫�ח�Q�����0�^(u�2���3FX8�tS������.�qQ\��a1���Ҩ�s���$V��(��n���w�C��]����w=�5/����t��_��Ke�N"�#g\7>/�sBK����e�X�slo��Z*�.m���$�k#�-B��Es,���W�W��y�h������'���ۯ�s��(���r�i�VtPm��h��zN�Йb�:�5�0,�&_�8��6�����uC�X�l8�'Q��D�=I2o�W
 Ŷu:y����UY� �i?��*���"B�u��Q���U�.BY�A��p��nZ=)��x��Х���!�r�^��T�*���������P���K5`�vE8 ��Z�;5~BX�CO$��*�e�ē�ŬWΣ�f%l�NA�ɀ{�#ݛ���_N��ò|�t��E�0椸�]9��W���X¥�#w���8����a�I\���.��"H<9�o��J��)��4���2�(�+��_��d�&t|�eZ	��.�H,f*��`ԝo��W�̰ERE���I�;s
 ~��_tm�R��B��RC�I���e�6I[F>�.������qWXm�����	�kU��	�TB8U��_<t6�0���^�k���M�KEj$���VY��`��k"�.���bE%#�<0ޞ���_{�ߦ�V��b�DJ3e�XB *�2���,{&0RI���Լ\4ο�>��U$D#��/�W��6���éº�3Yc%=&"�o&wb��"��ȇ�HW�Uݱ�+�L;�{y)����(���X��a�H����ZO_�_�Y�utfB����x��u�=q���C&�����Je�4LU���Ȧ}�$��j����NC�.&^��l�gҮ�CUHH�A#��Y4���g&}B�ޑ�S�\� n�]���dgW}�]��)Z�1$Fi(������W�����l #���a�1�,jUL:��x�ﾞV���E^I���O���u�E�i�f}&jy��΢mMD�݊QX �k�+��p������Ċ�34_����������]0뻣b�Y�M��(���5q:����_��>�J�e�e�e\K�3���]����GQ�s��0��p������uyy�;v�304�
�`�q�2��7��I���9��՞E�@p*���4<GkZv�E	��d�_�y�	r�����k~�5�[>�Tq�Ft�ד�d��JN���-�j������OVMߠ�sf#� ��ƽA�/&��	����;�e�1�<=��Њ���HQH@�@q�5���.#� 0�u)HA2�,B��>:���X㊎3�X�nopff�R�®��ւ���[���[��0䜥Yٷ�=�d�~�<��Z��Uրc��lK�n�w�q���}�'��f��y��Q���N���8`��E�䚊{���^��d�H)|4��V�220:�q_PG�ffY)N�>9�d�[%�E��k�{�mz��?�ψrͫ.w�������nX���2���P:��y��B�u/5V��%l+	ms�R�G��w�:�1W����/Ž� �慞޼��0��b�F������6Ș#�wJD�LY#vX����=�^�R��av�G�G�&%s��令�$]��"�!Z$95�7�I!�����r���o��jA��u:vn v� �v��=-`�5E��U\�$)�sV=! �G��Y^��U��3G�R�G���9$��Li����Vƴ���_�7�����^-�8��|Z�%�S�t|�*UX48��b�Z�ݮ�d�|v�o�ɯ�^�+.�r�L^M\F���i5)ޮ̇�iߴ�|f�H �v�	������a�?Kw�4�D�Xs��k��<�S1(����w,�b��R��&P5�ߒ��_A����Pt�]�џ#�|�a���N��4|T6���Br��9�sL.�LkЃtiݞ�ϛx��+ab�5/��G١Q���ph���q�^;
~��m�U�R_T�P�T(m���_g:��y}�j��N^���9�uJ��H��32�o�}%m��IjQ��=H�1�J�?I��2��/AI+O��f4�-�B�w,qǨ���-����I�#^"�!m�K-ߨ8��T�N|kH�n�AD9�PL5l�6E��� )S�3�\�]4��*qR�G����[O�:� ��Bw:��6W ��<�kl6���A �]�IC������(�eĲ��)v �IAf��m�]C�"�ğ���9[�a��V�1-q����(?N9�
Һ�xR&b$y�%#3�ɰa7�V/�"
�t�����1m���*��>O��o����sx�܄��!���@�5\���@k7I���ݾ n���y�I���)�������d�_`�	����6�"�O\m�m�(Î���3<xso�4�c?�����Lb˒����BI��mNfp[���#�!z+��OfL���}h�ɵ�WY%84��w-���'%L��$��+���hz���� �RE��P-@8ŧv��͜��1�ӷ�	m�6q��/5����|NsC�J]Ȓ6ļ��dO�ֆ*���냚��%�Z��i5��Kόe<�1��<��[�����ߛ�,Y�>����Bo=Uy��"sm)�)D�� "˄���~XЦ���J:b퐳��%��elMn[t�9B�X�o�	~�J<���4��/١��6�Q��},���J����[T����8R�&SJo�W�~��ȸ3��=�K.�_k�2>��Z�)֗���\�7y�p�Z�k��}�d�8�%�4*ٵw`{�����F%M�<�饚|2�q����G���v�����~�0'.h�[^&��ΪY��!M+���������0CZ pp>�7�V�x�� � ��U~4p+�s�=�g ���q�D�c��ڧK�`��崝J���G
q6��j��((��a���?U��GE�X.=97_�?�v���6��yHk�����S�����_͙+�}��yߦ�FFڐ!N�Q�ǟ^���(�X��T1u	��<�'9�� ���5 �gٙ�U���M¯.�����D��v	���_�b��ďa+=�����.a�1X���!�>�	�g��h��6��rBB ������ڇ�l/���^��ݛ�R;XΥ	txb,P�����F�ԟN������;�b� |K��W ������N���f�"�*@ez��J��
[hs�V�z��"h�;�-��q�D@Kn(�`vp��.z&4\i�}��Զ�݆c���y�<Fi�V�C�٪�m`;�b_Ż��j �CvGg�R��Ŭ����F��ā!	�ޥcS��r3xǓ��fמz�d�-������4yjnIH_2⩎}���;݃L�_"��]D�m�$�|9�E�gg 9�Lu�� ~��?�r�X���u(��z�ӱ�a)���\^h9�PUD��T�R2]f8r�>��65�p��HH�c�x�"�5�N�{3p�*+�,�9|���=�!��2V�µ	u���ݚ��4�pJB�,��[�ܥ7	�N��ύ�mW����t��]�⤿��\:56���� zf��p��$��m䞍��c(Z!񳊔�ݲ⌲��� C=xl����l���4�}�s|8?�Nȋ���ܚ��GeH �^6�H�A��g&fL��I��M�?Q��	T6BT�����Gzd�sN���6�Sz�eHݙl��:��Ίd��ƽ �zQ����鍼��E5��H�T�vCg��t$��l�ѽ�i8�Ӵ�h���'Ќ���zb��4xE�n��w�-ez3`�>ά���R�*����P�#��$��Dq��L�=w����~ ��0�N���qv���g�1C�U���b�3WV�hK	����>�U���<�W:5�ۈ�J�_>KO~ W�@Ȇ�q���8�٧:A�����MB����8Zrr{��x�hQN���_"���;���O���^�j�����T�J:���s�
`��g�i�D3T�4�G4؉D��}�w�)mmU��+rU4�ē=p����,ekp��H���ǻ�*2}���C�͑S%Q`ޱXN�pCǪų����4C��e�SfiF��\�5�5r��D�SТHΉ�.��4�2�D��2�G'x]]"K�����E-*w4��|�+h3vW�07�Trt�ō�u���Q�r�����t�G�r�jƬ9;��S�/�=n@�O�����ӄxn�]���X��W��^�'�]�c� �wP�O1�����,�ʤk��� �c�����fq~��z-9��@#�䴍�NG�zIr��Bʄ�vȝ}@�j�I��䯊r/v����S����Hڪ�<h�u�1�pn��h��rO�l��N�ɼF��LeH�ؙ���+�4�D��¸a�m*�U��;7LG	�f�ed���,�a3)_���I�mψ"�TE���<w�:m�PeB�� �6ȏ�Z�r2�{T�o��0(P7{*|�v#�O�	�V���jmt���f8?J�� ��r�(�����E(�֮���l��4���q&y��<{���@�2,JH�6j��T��"��"ױ�t�3M���V��Z��{R��G��=KT���}�nұ�������Z�<��~������P����eA����I��e&s<:}35lh;t�z4j(;w;���UC�)ѣ�.@�iv0d�p�a�TUZD���ѓu|�����JC�i]���3P`]�༠*�3�ɧAoزI�Z�V�b��lq8�o�n㹃Պu�ñ\�N9�RF�zbŻR+�9h���oa����N����V�G��k�q��o�\�3���o���@����]qd����_ԫ��
z��xG�H4�Hg<7F�%��xd8X�&�8@e�D�)%l�m���(F�������3�S�tʅ�x�4�9]!�њ&���:�S��h�)]=��W��Wo��]�{Ğ&lI������n�84 �r)޲�S&����B?_=�o���Oh����P��B,�+���Q��[y��ey�n$��ju4�8}鍥ޤJ�|DĹM��ȱ�1�Y�<�� z��G\dOA NHZVC�n�A�ß#V�� 5�W����<5��g5�2w�%$��-�Q�Ӓ��PBUu0R��C*��j%kp;ɡQ����n����0�<ˉ�ϴ3����n��q,٥�Os��h��x��'�J{k
!����/v9q������-�GO&�p���A� \���Yu`�%u� �М%�QKFx�,��^�BH߂�����U�g�O���[h֪k]؋����^��c�16��RP��K����c��ΆvP��1�-J��Cl��P���	�3�U���
L�G��X��Ä=�r�@�u���t4jL��%���\]�v�����	����+�BL����)%G�=!c�G�=]�F'v�$����=�$��e=���H�d���̌����,�ݷ�{��(���f<M^�2	�ϛ=��f�������x�D�[x��CFvs�,���\hB����1�~�	�z�����6�JB��%OyZ�����"�S��\�jm�bMo�f��9��4���"oЍ#D�[(0�6i���~������ �n��`~�á��������&$a7��Jm��@n�Y�X"U�L�����F�N����/!�`ħ#R��O��k���e�J1@F>���S����pt5	�ohؗ]�H�0:�_&��`Ny� �����gC�E�Qܚk��Ԝ[��h�!y~l���F�#�B��
"ԛ>jspyP/nAɹD��B�37ހbƢ�4�Y��5���(�g vU�������lut�������`�ً��6G��B�+��ߠQr�f1bq����c)���{�}v�L��I� F��)j�(��F=�hb��;Q]��ǹ*8�|��c��\�pY0DZMf�} ۑ�;�}�� ?T�JO���W�Ê�B=���'�g����K:��P�`
^��9r������d޽y�:�o�g�� C�&V,0�`��I<
�^��7�*n1޴Z#ŉ؅δeTO��r����5�BsIg�l��k�](>�^�9ɀX :��O��}��܊�3��3��(J�<;�
�`M�ӌ�</51�-;Ieb$G�Sh�A��9_�$I< �ؖT�w�Q-GQ�@*(��;��/�6K�zq�d������OPq�,�7a+[~�ko��k02"��v �5�ē��)���Td�N�(�F�N���;`�knw�B�������+����wp�we�Y�!��{t����ǰܼ�;��q��$ÊH�f����S�%g��`C������E�B-��*ې�s�M�]V��L[�t�|��d��<�%�����7�t [�vΛ�Ao�a����"=�����v�K�W)F�n��
.�B":)RN�e9�VxX%3؈��J�c��I����yB���١�6�����<=Y ����]Y+�=��8�r˾z�+����?-�EM�����^c�+Wy�ֵ�)��� ��C0�!S�1�e�Er���΄<{�p[*��/y
��T䍍�ǃݓh	��?�*1��W����������/��ID���+�ʆ�?���S�}��`�H$ilC1E�{R��.'Z��/<9��W|x�yV�Va���}�)�:Ȗ,���v9��������Y�1�Co~F�{�;�	n���N�v!�!?��0|��ހslk!O��l:Hv��f��Wc�:���gEع���0�i��'e�B�+����0^��@ @	�ByE�
��������QF����G��ڹ&�4�PҀ4~�߷G�4�i�Ik���-�i��e6�t�	]�!�B�f����~�B=��yF�,��ul��P�I���u�!�1���\�$�t�6-���<���9�Lf����rg]��%���JD��}�����BP��ǕY���wf]��hU�ze=�=ה(E���~�0Amr���zR���U�����w�_��+�p�b�����rCޟur�)2���BY�V�0�0�F�e'�a��y��L��R��C=��E����9�+��M���y1���$,���W!�l��I-T���^]��+T'�Z/[��&���7!px:����&U·�SXo���Z�S�B�Q+y;uKp�<d_'�*�AT��^�n7���m��I^JO�����y*M�98QMO���D�	��6����&���WU'p��+�jC׵W\O�%���ԧ�M�gL�Z�Yd+�w"��'�[NTn�i<�U�@g�$���B�|��r�%%�f3tO�e�dyCMY�l�Y.ҫ��JsYC��d$,�������rɶ9ś�lsH.<ܣJ�IVa��'&J�w0���)2dzjLb=���������a���&��O�s(Ǖ_n|���BC����`�q�9�R�/��T",b��n��0Qkzڲ��6��L��}s��v�Ó���W9pEm�N]��w�Ö5*:넠��g��q���¬��|Rۯ����'��l���g ��Z����0��hJ��x�;#k����Ļ�C�p�l�\q�m���3�敳�!rƬ	O`-��\�$�<gʇE���V泟�B^I6s������8�[/�K�E��LQ��w1��&�b
�'�����E�m����u������M\"�,�`P{z��#k�v�}w�!��[!��j��-�/�@w���(E�}���I����	ڱ�w��֒��39@Og�`zju�dΩ��w�X)I^� �hǻ/_�1���B�����l�+y_hV)[����c�k�ڛg'�w{6F�(gɭ�Tğ�����"m�k��f�/�n{�&°��!X�D��H�U�vRo��|/(�#4k�HO��(��Y&2�U9f�L�7��Rq�L��޻�Pw<��K>�CoX_`�5|'X�~V�nR��פ����u������S�@�p CC�x"��ȶ�t����.�wi�	��z�9P8P*ip�r;��-�I�,���sz��$�:��̂�XZ-����i���C�S5�v_B���b������d� �Y*�I��~k�֘��W��;��褁��@S��Cʼn;r��B��
�*X��GPȺ���V�L�"�韢��<����Yۊ@�Ml�'��F\��7���j6ޝ4�aJc��UIs�M>^�0��B�4��zN���r���C�%W���{�ʉ&x�����#�Ly9A5Z5�p �aj5���e�)��_ŏ�Dv�܍*Ы�n-$B5���a���@��_���?=m;w����V�v��B��z��"�ܸqF��4�f�d�K�.�+�uR�Drt'z�5�5@�T���-D�?�d��a�B�َ�gkZ"^E��B��""\&�`UK���P���ZX0m���qm�?8�M��b�JtO�������Eݴ��p��rӉ�єE=n����Ś��b� ��!ܺl�	�n"](Q�C��]������]��Ӵ�āDF�1߉�.���+��{Ϭ���8�+��Eۚ.`���l��ߛs� b"�z蘆W;��ɲO�0*��:�Q��NNg{��Lo��t7�9�
q�#Ԟ1����n��^D�rHdRv����vlK>wW�;߿B~�`p�-W�؜*I�q�7�N����4���[k~��~W�y7�E�ʼ�JT��J�ŋ�R��P�ai��mAcVKW�'?vʊ�Wd����1w���b>�R�>{i�<Չ�a�{�#� �O��1�<���X�Mnp�ܡ��
���b�-���n0�dS�U6M鳡f��bA$���L��wQ0��;{���%���k�s��^]��49�5?�z���H��ȅ��0��ٕO����ɞ?|v�B2�u-��R�K΂���4�X��$bu�	$:l�߅=[i����@+y�;u��f/��<���³� y.�^c[�/�I���P6����)�X_72R�j���B�^�eN[ߦ���Cw�1Z���mg2W�P�~���W��񋁵v��gq��r"$��P�.��j�V���צ��[�%��?D�Mw�e��]��>Qۙn�C%�Y�b�H�`�G_�Q�����:c�b�a+�8�K�	�Re�݁R���{��E��2*'�o��SZ쇖6퇘*�P{���9U���wKr���E�eO!֠�]:4T_�z&�?�M�� ?%dݚ?o�����{~%�KD�7�IY!�A)Olv�������H��@f�[���B�K�H��ݐ3%�	���Cy8�[�K͛
D��^�0u�棦"+�����%�nV�r���d�52<�V�#�>����&+��E,Ub,�@�.BGA}�,���� �Ak��il�V,��Ｖ*�1U�ёN�8�r��s��	����8��<0>��S9�jhe���]��N��h��xs#�����E��.��O{[?�{�3#󂞛1�Z}ޏI������ʹ�6!ݛsdX�Y,�5Xx���rG����=
Ԭ(�TR�V������l���#�.@Ȇ�k��JӴ���=��09$���D¾+l��f_(.Lod=���qLwg;Ypk�I
�I������oU���Թ��l�������r/1#8D�q�4^wHn���A%�w=�"5)e��e��m`ou�d��I�R",��<O�������E����9Z0|��NW����Ԋ����L�=�\���b���x9�`�<W���	��AD���_F�Zch'����GCM6�6j���?|�,6���jg	�1���aK$�ON&�,e%s��Tw�p�"8��#�}�3���R�^�!�PTm}��fns�%���0��ž�xP,��ݰj�;CՂ��94���Y?rG��v���Ƿx�J$a't�Q��8��o�Ǧ��Uqܯ�j߱�z#wffO��^
�W�i�W\h��$&�X."p��+����$�͂�
�<���<�Kg���Wf��@�݋�`�e�9�=�mYB�βT��؀� *��*�B�Uʹ,=)m0�'똂ipp���J��)EǦ#�p�{��&i[���HS@��3X8�s�9��Bx�YҤT����(��^�]��H{-����)n��yw���S��kf��4��_"U2�q���r���bZ��!Y2��gE�M���x��a��P�_�a��0��,M�$�-h��T2�oىE�
��_����E��۫ �?�#*��-6#��:�ό��^mo�p��C���a\���ē�ʰb�O;�]��CIz��'̉��=�����d;bN.n�kF�>YY���:9ږ6�E�1ϵ�
č�W͠���_�8r����������_r{�����#�L� ����f����B���d����R���#�q�N%M��9�ѐ{Y	��9P�/v6��B��Tۀ�FdsrW�(>�cx,O�zݞ�X'Z<��W���
�.�8l��=�R�cG9;��6�ħ(�${���v�ft�b�
� �nFy�
��������J�T��1I��1\�M�AW�i^'�GVw���{$,J �?opl��T��e;@��Z̈́��g�|�0��]���T���y����e.8�ԌZC�M��xKb�WA��hBI�(��ˁ<�h��#����ZL�z�����+��u_}
�#���d�k~$�C8�<(?}P���>��Z-Y3� ��� ��ѺN� Dae�����+�1�^�#����F��hX-o!K��u�Գ�U���H��!.ĨNfZ�A^�׃V�ë6oD6���a����+<��OXQ����'�{s��`\ث�!�n#[�X�!�#�pF�ӠS�:�H�qBlq���.L��_Ԫ��,%��Զ!j��hl�����RM��nu�}��"��I��SM{�O���W��?��n#������q�x�����sAIՑ�������ƅ�3;�x��r�I,t�M�_�o�ڢ;U��v�	bW�9���i�2I|�싯��AӮ�>��E���"�V�ǉ_�Ӣ�]��!5j`�\:�s�^Y"�H�QkY�i���Vy����+O3�a?�p�&!�J@e�%�t\E<R9��������m��e�_1;ߑHg�Y+�"���c�![��
�B`Q+�4�g���p0~��P��< �ݖ	�z�B�-	J_�R:@�*k�B:��:�|�V�����>	f��׸�����n�\���况NǴ9����t=���]����_0[U"�L���b���9(D�]�
p�����1��?����7�����������'00������W]`���紹�$���pf�.���p?^�!/!o���qf+%��f�B^�Bq�g��Xc���6�=�z�)��)�u`�i�0��Ӏ�[�Ũn���p!:]L�K�ar*��6�b}�.�>�#ૅ����(o��.�yz�$�3��D_Հ�_�X�uP�rݥ�d5��a��<��5؅F���<��0H���j(a���r	w�|G15��N�	_7�A���٘�;C�4�#�|���O����X���2�o)F��n���j������������_�H]9T�,���^+ҳ��=�� �s�R�!�y��d�IoO��L�s�����;U�S1�`�5g*8�X_����h��Rrx�kl��6��$��N���� `�偏V;xEFX��a A�����\�	��0����5A��)&��PK�Qу3���[���F��OY�W@�9w���9�i��?{4FO<׀�"�^B�����f��.]U�/�����P�a�n��nɹ��+Kw��k�
zR)^��w�vs�����m�V���v��O�E�w�E_��#4�B@�i��S�y�'�L2���{Q8�����5k}�lb�۴�<��������z�i����O�풓��	��d�Z7�	C�֡	q�6Y���r��_|H ��hR"�W!��m�m���R��o��b�2�Kz��$�b�}�AgW�,�Thf����4�E��3gR.�Jx�MC��i�>i��d�����}���I��� ��wE撉bP���N��7���d�E�6g^H����lg{�ݍx��eA"�~���!�H@A��"#C�;~���X�9ۼ<f?�P�����U��0�q�,��֎r�W=}E�&<f��B��WT�`Ə��r���ڝО�)3g,�+��џ��-N):�g��?v<^\�i���WQ���Y����_�%����n	����X��H��n�Wqi��+��9(����6�n�!��m����J����*9i���3��;��p��$���V����bp>%�K%lJ�+g��yQ=ۤΖ�LE�-R�B�ƾI�M�$
�d�B�ڿ�@/W���{
V���9��vg�o�DH��B��� s�9�Q��}��Vm^�͜�l�8�ZiމO���gT\��;ʤ����:��"���%nl���{E��rϾ G�l�@�GB_4����$Mu��#HJ�������i]����N��w�t�ݛ�G3�z2|�_vˆ�=���S�M���%���@U'=�Wۦ���y�U�3 )��QBŬ1������������/#/��A����ϰ/@Z�~^��=U=.Or�IދJ�e`N����R}e�<����'}�.�L4��4���~I����rK*a�g}�����7m��&r,{]�fJ���z0^NgM����i��y���Sd�(�Dkɬ�`������mb2bzd4� ��kb:׷D��px�CBEG�Կ����J�joo�&1�6��ey��S6���ѧ�@į�2)~�J����p�������E"Kߝ�V<]��l1�j��q�#�N���gR�N�V���c�$��se�A�j	�'�\�<�{^߯�x�p��h]����ח
�2�x9�Z^l��PJ�ݭ-!�|G7�#er�*M�'�6����W�M�ҏ��s7�'�
�����|9>���d��!+� ���H�k�p��eq�ᩔ��i�X����$��yВ
�d��8�J��!�7ύ�s��Zn�SmQ��[��ڃ�u��U��ͨ�G9�&$�%��We��u�%�K:#��C�4�W��k�mL��i��Y�9a,�����HfшI�x�c6�Y�}o�p�#������?��Z��l)gK)�Nu��<�b���H(`>�q��7`��7,W�ƠQA�b�G"�?���*�'�H�p���# ���O��e+U<w/�a{���A9Iۼ>�� g�6$v�� c? ��@�p�Rxt��.�{&��*�*�JV"�֜}�a�y�n�"T��dS�W0ꦛ�7�3�]m-	y_�0�Yd!������hG%��,9m�W�6��E����C	�[���$}q�ܯY#�,���Z	�~�s^�a-�4�P$^�ft���%��wr����,r�C�a�ic`[fǓP�7�����KօD�ŴŦ�O�MW��ƅn���c��zGs�MXsZ�Kv5:h9��Qh��N"�I�9%�� l	�M�WՏNx��_��L_t��z�֖�ۤ��>��z�Z�'���C!!���5�����*f�W�ԫ���ײ��F(fԕ���<����LjMH4���f�-E��� vT&�݂;p$��0h��辻F���N�
w��]�v��Й�[D!Z���9 �h�h��
}b��93c��ZX�.�����6����O�H�b��������Ή��-����*�T?R؎zU�����:^ט��:s�D:��P�۸{�߆����'
'��C�<�ֿ]q��t����Ɠ��hR����O�1���&	�E
�z��n�+���������0����f،��I�	e�|G@�ɜ�t`zwי����m.n�~�;��K����q$ͻ�.�YN��:�E�t	��Q82�0��mq��G�`���h����]h`_�C�������C��n��o%�M�e-�Od*��6�H���j��'婶'H��}�Ԅ�t"F>ݢrEy,�M�#Sx���_ф�ie�2�	����F5�
�H�B���EoqS�(
�QQ�4Lہ9/�?����=�Ea��]�����J����K����MN�2{����N�
��H��ϑ�	^/r�@P��;	�}����R
E��e��N
���o�i�Vg_E�U���U�aq�4�wױ�X�R�,h�N�p��?9\8�s�����ʞ����rס���}����m��O�G�I���[��W�5�l\y-M~��.Y,�>��Ќ�Z�'cW����^
���R����"��^�b����:ְ�,f>.v �p)��]S�D�u���?N��`�������Ԫ�xx��-�>���'(xO���[E���W���P���HC�����G���w/<3r�Cʧ�ùO��J`_�%���~���@���_e4�Z�>��Q@^?"������S?��(�a�w+�;3^�ƿW�f����T�vڊ#��m���5Q�3�Xk�UP���>��j�S�am3i�Ԋ��H�����%v��Jy#�=Cc�g*���Ȅm{E/����lk.ʤ�&N+O�e��xԨ�u��D�@�T�oj�60�Q���}`f�~E[���r��0�:�4���;=�S��Ʈo�<�o���1cY__=�L��M��ʫ�߫��1�J���u�G� T��.}!3/d2�I�?5�s��-��\��C-4� )�4(_�;�Q�X�[Ђ$X�v_���0�3t��ޫp��_It�:�k�vrQ���d)܃Z���Eр#&6C�P���\�̛��,X��X&�1�9��� ��laQ�f��(V��%��Q�p���{3���"Ib!���	�������H��X5�ھj*�����WQ�����@�C�x�N@W.iP$rx�#����~lC�v����%��BG�h^����B�F���d}]�5#��kvςF����y>&�������w)97��1[�z��z����z��Y�h;6��+PL	���)�3��LN�Ѕ*��P(���7���B{oN5yvՐ�\7���'�N�8�$+x1*\��K����R��>��O�^Nh���&�r��#��n�7��S/�O�J_01t�����fi�J��?[5� �:��~��R�Ұ΃a�vMd�Ϲ�\j(#:��Q���/�C�����*G��g(_K��,\XS
�qԁ���oY6�ʛ`nJ�h�;HNYS�y/�I5�3�-�������~$[�(�#-0�[B=��Dm�r�A:C�y>�����׃�|�B�����q{I�H�TW3:���b駅vɘ N�:�d���~YU�yq+���lכ�4Eز+���(��l����>"��X4�V�Ǐ��{�:�ٌxb)��[��k�$���Ucp�	�8��KՐ��J�$:a����W����V,��.d<�C�����7�h�lh9��)VWM��>�L���Y���x]0?�L�����3�����Iz1qy�g�#NKt���~�UZ�^�D��`zN[,�>�ti�Q��<���㗫�JH�i>����zl0!�tU4wQ=�e��9�<�P����nn"�29���`�I�y�q��&�4�4~��@~�� ���*�v�kDH2SF��p��:~�f�\���w��w����2���x����Q1�#K�Y�=��OHi�M�������ʰc����:6���bz�,��!�s��p�)��1�ܰ?���N����6׳C���v�ej�͗z҄�
(�mI�Y��9�gU|R֘Vp��mWk�J��F�����Z�����S��$����s	�i<��G�Z�1���%@��l�����Ѓ�y��˫����'���
�+��ȏ%qRQ~�"4��;��p�x����/A��e���J`���	[5��h��C֩k]��ȹ��#2+mš ��^�����Φ R͞�y~��fsq�Yש[���-�vB`�1�����A�S<}�&�Y���(Kޏw4�PS�Z}�uJ��g��"�~Ү[]�V/%���\�DgD��$SY|]��ztƴ+ԓc<�S�4��\a�rz�3߬@��ͷw����O�1a�[���l���]Z���57��v�Pńf6TOa���<n���^�z�e �����>1*u��S�]#�`ݳ��mBr%Ձ�ҝ���!���y�xԜp�B�ܢ>v����}v��Üx}rݰ7�����4
A�;���|3�_a�>�����t>t�%^%A��()�j�.�
ek�4'�D�!��%~���qX�sg��N8o��*��T:NA.a�k�O|��H��RiP�O�hp��6 �S/^�M�(]�ԇ��PP����jT6.z��S��MƁ�ϊ��n^@ܣ�C���x.�����*3���n/�VP���o��H����))�2"GK�"a�wD�4Cy�Y����V�5�G��[6��nc���*��8���{M��e���t+�.�Z����1,���$�S"��b���v�XW�1������F}�KO¤;vN�Ym1���{��yEV��"/i�.Ԟ��R�BW0��}���6�77/��%��y%���E��I��k�!����J�=��[�+Z��`�˸�i��y�)���N��M��~����:Xژ���A���"�@�L�Hҷ��@hm�J/����`��l���|�m���S����ž�ፘ"ˤV����so
����!7�5�L^��Q���U;/cI4�����)�!ai1l�S�%4M����ҡ�~�m���W-/aAҒ�/lp&��?d��$_��O�(k�n�T���-�8t��n��W�I��iB�J��!�,�S�S2�џ-��QL�[#��W7��=��U&N���U4n�Y�q�2ӗ�6�9���KX�ɷ��	l���X+��h���`D�8�J���9[zla����B&���ܤ�A�3��`��($��P�t� c�h.��yZw��s�x�����l�}L��q��~N*y�9�<���Ş�-By���)���4�ݡ�l
�I��6�w���
j�q5����XIfϚ�G!���^�>�d	jgK�뇫jv��H�(!�kjy�UL��Ò�k�����v!9�2R��̘w�w�!CoN�Z|p̩����<!�s�x
l>[�A�ht������9��P�pD3��n3�x�
)��/����!}؏�ϞH2%���)?�D��^Nu�n�4K�u�.�K�]��;	ᰱ8 r��J�ܚ��'@�.���Cɇ�"&�/�wq�ZDP��V7�����?j�PA��v@I�b��F�jMk2�=W:�A��TB|�ۨ��Bq��������S��ς�P� Ze�WB�� �?�9דA�b��W�(�6Q5�6e+���=�1��ŰN/?�m�I��ݳ����+��!\3<,���S�A5��&-�����?�T�$�����/�!/��{a!]���Q�8��'<��5�뱥�eG)���(��٣{n��n:�fgR�0޹���2��}n<��_c�B'V?t(j��->fc�BeP���o^<(8���nǥ��Wæ��,f�	��<�X�8B���̆�Ȍ�7SH���Ы����IvͲ��ߠ��w?��&���jw�a8��U��q�&�ñ�Z¨{�/;�cC����b��4�Ad��L�ŀ�'q'B0�]e��}�62�A��W<����rj.&x����������phḄ�b�>���P?���=� 0��+3/�a����oL��K��H˩_m��RފU�!�H#E�L��:�4Ξ������3�e�nK�ZX6't��3��߁�W�t��{}ٝr�����SM�U�<�`b�X��f\��N>����K��j��f$}��&��蔪YU]ŵ_+��L%pIa����) �ۿ[��s$�!���L�̀;Y�7�t��V�(�e�V�;<������0d�@'\Ά�9P�i��3�h�N�H�s�P�Zl�y�tD߾M�e7��K/� �'��fuDD����;y#˓b0�Kgl�
ى�e��~:�~�[A����9�]!Z��<C�,�r}��MhH�	�|)��(�4�$��3VSl�<���[�t���9b�륽'�'��S������)Q�����'=
N~D9;��#��*��xs���l訛l��k� (�_6j�X�X���Q��� �)4�0�k9�z��
�i�|B��Z�3���ou޹�Q>#Jȭ{Z��7�d�4n	A�S�-�MkbR�Иf˦<�C�!��(Q�ƹ	��N��K'�U�/��p�k���E���^[9�4?�����bE���"�G׵ $JT��Z}�DkPki^qum
ZA��2��a*���I�ڃ���x��7��x������c�OX�x�e��,!�N�F��aV���%(8oR��4J(	�.%�Z}Mq�]��烞�	��3hI��ɷ.��uM�q�T7��~�P���3>I�Yz� �	�}��0��2h�5O�a�bB�?&����p�*�Ġ:R����A#7�˼Ogک�kc�dM�v�:��"(l*�,.\�����}�4g}�+�>�& <����;�2��ҏ�2��J�^��q�!<�+�?����?���h%�s�Z5�rE��X0��g�����Ԙ�U�ZP��9��v]*Z^d����]�,byV2��Q�j��>J~y��|��c�4WP�Ocbv"�,}��i��;n�;Ư�Ѵ�h~�da�y�10dI�a)13]ILY !Zp�'�k�1�Q�5�w%��Tqϋ-�!]�ق~҇�q�q��x>dnf2j�j��}���H�=4>�����4�݃ o�$��3��|�c�o�=�v��x6��i $�������r� �D��J����N��t�[�Z�	�����cwA��dk��"p��O�Q�+ߊ�KQաG�?�e�ko�o�A�(��N����)�/~p�'�x�]���騐�ܨ$tk�Չ�KM����K��ؚ	�'���N���5��G��wq���S�h�ɷ)�^���n�/K�⬦�ȾÁ�V��:���5��p�Qe��s�	O�򐋨�6��a��R'==�,�%7��@��A8�_���/�	��:/W�$�p�V5�db�!5A��*��e�.�����e|�RW�V�*!Gj�*�@�e4�A��vj}H�|~#MCܲE�����b���8Ke=s)7"��������kG���z��xy�����tVk��/{e�|��t~7�f��k��K���d���ľ���s���ݨK��
|���_����ڊ�#� ߀-Nmq���p��:mAf�" ��(;����-H@�`�U�(�C��cпD�ϳ�78Om�+���VD��;�(�C�����Q-��s����5dz�K��
��Z�*垲��{A��b�����y8���Loa����[�<W�D�����jgYm�4�1�ZS�[3Щ�v�
��%l�'
=��p��_~�~Wa��N����dʣ�_�����s�5��[���{�^f��E��:m��Pa[�o�*�����e��Ş�f��Yg��,:�J .ףy�ɏ�ǀ;��$B�� O����jO�"�_�d�pu,��&X�hy��3�b�џIM��!�����6!(�w9�b8〧y��(ܐ%�wCM|�$7sK�?TF6�c�e��%�������AR�5~}�u����K��v1a���f��$!��6�0�Jh.���Ao$��]ކ�kt���24`)
c����5cW�)��cWH �ܚ�����F�_T���t��?h�!�+���@��W5����ηٯ���"Vݠ�]��H��T�oN�x֡|0թdR>��$��4��X�@���Z����*�wi߄^��Dk�%y�Ib�8} 녇�K��W�7e��q�8g����k�ĩ��!,����L�2~?b�S��[%o��3A��㭮��WN���-���aW����?y١���j�3A��)���N�	��3���;�:zn�d2Ri�*z�Pi��B�e�"��S�v�������-�(�����/�6l�8�|��8�������S?q0�M�a�� �ƻ����%IO�b���]�B6�a�e�ù�Z4��Gs���虉[���ҘK�ҵT��A� ;�^Ƶz􇑫����-�k�'��GhԸ܏t�����]/Rllq���gִ�r���F�j����t�g�j �P�~����]ԥ$�2Hh�Yn��;��d;�b���ɝf��:\�u��j"yO���I�e�I�f�|�l�Y����J�vSQK�S�+ֵ�~��R��wvD�c��_R�&��B}z�9JJ�]_1�R��t����,n���]4Y>�)vO3 �MO;|��\"K{-�)Ӡ���P���g��PJs��4����s�-F���cD|�2�=�UB��.����t�7�|:#�����$���?��AZh��*d�<{�����٠���|�����7LFB�9K�]督��o�ռ��͐�.���/EM[h;�ElW]z��W�!*��b��BUGr�=.�C�j�N���4�n�u�n�T�Qt�����%��� �hx�#���R�o�}y�b���ƛ���f9��b��}e�_3�yHl8��<��+��u:��B�/�E���.b[�o�f	�י�7�-#�_���P�r�9���^ 0p����)��}��/�?h�(JZl�#�4�������ո;T�|����lmX.��i%�K�Sn|�M!T�i�%��>�2	�Qn��1��`XZr�Iq7Pa�ipF���&�Q$����b��0�>E��n]Ri��{R�[��lf�-+	 3i��!���np�P��b��،���1���|�xWƝ�s7FG�8�|�/���N{T��#s�����9M>[ ��ZF��(^= ,��1뢊]4�͟]��G�
��Aƃ��ǖm���$PU�F��ke+��w߬���Z\˹��*�'N ��;�7��`+��"�bըϸv9��l��	�;g��3
-�5Z�a/�V*w�$r˳X0�q�@"� E�k���������g^y"��U��(�7��g��me���3a6�~@�7I˹�i)���rsLSA�4��ՃCr�M13�!�eSth'�=�3���yC���fx��!�M>��K^GL�$N�� ���Z��_xi�b ��Lĩwk� ���˽�-Q9&��(���w��歽�%'z���Zrt��0^˥��"�As�2@�C`	�TEc�Je��Z����QӇ��Q��j�W�vyx4b�����H<��$��z$RV���`#l(������.`i�< �=��k�fF��L�}��<�08��K"L�PTG�����8��Z(���W(?��?"�Kۺ�R�V>_4y�5����>쇷�}Hjb�j����<��%�=4�E�?���ߌ6�p�
��z0�$�*��ql�����ٚu��ɒ�-j��=�r�*�
&�,_���ƃd���|e�_�XVVuchY��*���k��)M�3�"������`� i��3C�H��,��5�³�CQޟ�lb�a�PjqUQwZ��f�	��=}\�����v:�k�	��N��V׋���*�*�]��k��h�'�}Y�O]���<47�;i��'�J��q�+1�ʃ���|���u�/����5�GvWN��?S�s�����Vi�'��P���}�� }�)�
��0X�q��J��%z%��r�r[;�8 �r�]P��oc�(O���/TsԕV�:��,�����D�[#�C���w'lrj�g3���'>:l}�[gs�F��2l�|G�I)��_��Ĥ����K�#��t*@*�d�N!d<35е)���>
�2z������*Z{�,�Gl࿱q��e�?�R�$��E�ߌ�\sڹy�쳮L.{���X��E�=�(���'��W�e��=�n�	͞?*��$S�圥(�{�~��������^��W�ԧH0:*{��.7{�Q���ڊ�C�,�'�;�������Gэ�ON17��$=�y��p�/!��E¼���DE�� �r7����?5��B�����K4|�i��� ��Q��ۊ �uxt���h�՛G,9v5d��xb��@����_���Z	=!��Y	vB�Yi���1ȗ�*=��O��]8��E�/�W�Vo����dX(�*�v�O��p��d�"��S.��p���T�b�HU�Y��UWv���!)q�<As��E,_B��a����kÔ�iSP'��D+�0#�Q0�\� �@	��n����)�y��آ��o��po�����T�� ʺtBw�6Ncq���<W�K���+BH�iLquE@���V#ˀx7 �U-�PA0���~�����%�ЎGxJ�$��I�M���5�k>�G�{<N���L������OL��i��Jju���%2�c�3Ql����3)�.х���n���ǌyc�w�������S[�, I�hK�}@��`��OBhdZQ�
��W��O�s���v��Va�!��9�����R�7IU��ڗ�Q&�(�v���6I�f�n��|rZq��;��rW}���"KR/X=v�y��K	'P=��~�9caƥg5<��C)(Zy��gT��WvTPu���D�Kڥ���2ɢ��*�9�՚`VU������}U?I��v�"�D"��:c��:��S���K!���f���T|���%�m�~�HYkk'��4<��������s�
�6�S�f�|Q4�ޚ�����87ty����q&��Y�c��s�d�n��jJ;�Ә�ĲE��W�!�@��%�*B��g	-OS���5i��+�:̎��ZmZ��h:�P,�E}�"����Cl� !���������s�@F�:+¼��b/��#��D�#��ޮ���Ua��CnOr��5�T�؅��u����K�SP,�	�Pp&�~�M��b!b��rۖ:��&��8�\Ch�#bTd��
�մ���ދ��8���Z��?�g��s�N�zzM��Ft�ԋ��Ʀ�0}�Me �ObO��M8R����&��l�W�o�C5G��E/?qs�V;��ԑ�#@��U�#N/y!F g�WH������(X"��H�2e��!�Ы�L�V�����o�+�K<ă�s�U&�	&���g�?�s!����D�^��V���Fv
L��;
�3-�[C�[�F���r�>
�C=��}�)+f�8��Y��R���U�lYE?C����,�i���r+���S��;%+VD�������G��k��Y 3�Q.l�rGJn��(Ht�fdC�q���@�q#o�݊�ǿ��'P
m�r������=k�]��$j[��]�Z��=�B�!/�g��9fN�݉Lr{���$���(�^�ŀЩ/�tސ���=�ۊx�([,�껌��� S��M�r��K`۠9����Xii�����ׄP?�u�z5�W>�x>�`���s�K�������G�.�Wl�XF
[���X�&Ð.gG鯘>C*����e_�{�5,@��H�����{*�[ ���� ���W���%~{Fb����0RJ�5żeV9ƜG��>uV�I_R|��y)�M����I��X)���a)��چP�hy(,s����MgeL+J�~��.\X�/��8���!�c���i��L��j���}��� h��U�Id�n-79�2���\/�95�5q��?fAQPV{��Z��9�:�g<�}Swk)�K�o�F�6S�Z8ؑ�l:�h}MCS�����;D��] N�k;$|hί0�.�Xf�"�>ȕ��L�Te�̤��k�r�{r���!]�I'�պ�6�-F;0���M2�
lӠ���������Fu}�*2��tf�|�1E1���vR ���%���9���r0P0f�-��~�y����T�������������"�
�)�҄O~Wq�n&ۊQU`T�R���qȓ�۾-[���XF&>�ov�R�'H�q�(k�P"�@��GP+~<k�=�9�m�b����Q�z[���F�J�.&�3�i��T��6Ǟ�/��F�n�M��:��9���J8��҄��|eK��*�ckQ��`l�)�rAW0�Y?���Ӕ�X#�똰2�  i�3�b��K��\Y�2&��5��3)n�&f�8j�5s��sW(�o5��;�0܍l8��K ��~��W	؞	�Z�b�g�"�Z1�A��=���|�9 ���q�z��ˉ��>�xψ��2�	�p��e�=Ư6�_R66z��0��ľY���]��s��+���a����,]j��:�:����X5�<'&�d�'�I��Cd��ѝc�����J���n�Eހ���b�n1�a��-~����?2!P��?G}��EU��g�T����9���k��됖�<�	���cOȥSkm6���z�������k�$X�Z�rF��и�^"M�y��9˶8l��9��KW[m�o�5T**�
�|�G�Z(�9ύG��5h���j���w=�^.?�]���NS�oi���M�JT�j�o��)���k����ڍ�0H ��0
��5�Z,w����\����ؼ�����?�<2.���hr\��P�1j ��ۍn!��5�Ǌ�w��^uaH��G|���vJp��[`R�bY5�	Aya�P]���"����~~�v�s�����)���m�=n�w���9��N�;�k8��#-,p/K�?7���NKsܨ�ھ*������<�r#3�(�1	^������-�+fj���$j�WW�0���E?}T��� �K�	W�5?���y_�F[ĕ��*��6�j8߁LAEm�q%u���)o4��!��_M'��
�kTY���@���tb��&](Ӆ���;L�4Kj;�-��FQt2V�*�K.��,I��w/��XH���st ��AΜ���9�_��B��W���ĳ�����!S��e�!���k?wg�qX�A�p�5�Q]�T%p�D���_Ւ���M6g��qg�u� -�.?����x��o'�l?A�&���(@0���k���P|7�ŋV5@�&���ק��ۉ�����d/�r團�Qm0��y�=ǿ``c�O��+��&n�g*f�i��=��)�t�4�fz92�i�ȅJ�W��7d���-`&LF��1:U�٘���*/d?�[�-��������/��h�>/CA���<�A���m9��83F��/d�)�,���J�:m�q;�)i��`p�ꤔ�z����-ѱ���򉒞'��h;�<\m��!��و�+��� *B��&�_��c�8$w�>�@'_������5K���.��Fq��=ZLD�o���B�=�8癡b�k������v7h%��mى�ߔ1^���#���X�=ު��[?����y�iN�T�<�@�����L[��S��0 *�B�=���o�r���!\R�{^Ԧ�Qv�����A���jI��E&���:M�^4��