��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ`T�}�w7�ɴ��劂�����'�r]ju��$X�/v�A�P��|��u��}�5eT���ut#g �>�^�<�[G�:�6 �/d�6�k�~�*;n ����'�0.\����},|5�k0q$�8w�q"2l!�W{>;������\��|e#�l3�LIO��A���
WB�ۙ�^�3hjTOO"a��� �|A+�����Cu�}nq�&��\p�7D7�Moi���7u�D\���������+@�VW�O���u�f�+^ PԖ�;�J#܅�̀|�E��}i�Dʬ��U��]�ޝ� $p�C)I*���c���!��q�ʃ�o��jSlӔ���yE;z:��o,W@��=Ɛ�������y���iJ��@�.���?��.�~'�2�o ��ó=��������&2�$���> +���1���&�abc�@���b�D
�b�����Xu�1�i5ؾ���ߢ%j�����y�4ߗ���e�6��� ��E��3`\z԰d��2|
���͡����h�f��>|3?S�!3�^��4ZL�8PQݔ�.���e�����>��#W�i�]$ !tK֨x" �װ��OZ�/��������>�Kd
}�4VrÖ��2�Y�CJdCd��p��@�v
X�&" �^�j�~��a�����H0/mcXzm�\Xh�
�t����5�igw�I���:i�k�q��S��_�kJ҃��ًP��D�a���HJ�ʑ�)8�R�(*ҹ����j_�Z���[�Ժ"}l�fF���>wFZT�(�}*3I��U@�#�pk�g��(����X����X�����>���3gL�i��1����T"1��&AS#�r��1[��(��r�>���&us�Ѯ*}U��\����:��M�b%�j��1[�I���h�;d���Lʮ[~?�eo>@�7�{F@�֖v�4���eϠd�R������~��ؒ���P�|��Z�`%l�G<���4a�^^+GSu��%�r�&�aq�P��6cT�h�9T�:�U�5w�cQ^�/��0W��P,��� C���`̓��83�^���#��߀1����G{�+���Ń�jk2�
��+���r�;4�[�hq�~�!5��K]ɱ�����,-��:/U����=�����Kl���\��t����r1�}R��n��0��[�oq�y�9�OB�K�R=3��;wF�9�<I�d��J�i���A��N�W���
��������c�`<2�z"Ȝ���&#���C%��X4v�j��T�t+�F����,��m�>o����\c����M�ٲd���|���3>53�9^�jZ����HED"	
qɽO<�o�j�3�^��ąe*d;ӊ����I�S}+��B.� � ��YA#u�!�0�oS'���p9��y.��}w���K���12���R��|��t�)�+p��2��cɋ�'6B��Pt~���_w������J�V�����[|�G=��E텄����j+5�I���Q<F�r����]�D;W��}���Q@���|JE(��+t�xYzV��t�-M��\ߟ�>��K ��$��l����t Rӈ{�$�(�pFLL��m��I&0�U�}�1�������]�Y����{mc��������U��$k
47�I묒�U
��N$|xQ�%����;e��Z7Ԩ.Rxl��Y�A�3`R����Gև3�78.�Աu'4]��q���4t1k"7�Z���ME�f>nJ���g��Q�6�%j��+o)��k{�#k,�B�������[b_����Y��#�3 a@^�x�f_i�܊8�']���VJ��-�Ո��~XӃB���v5�k���g�*};l��F?�i����2�	E�6f�Uȁ S��7���/O!.���\�E��p�G��va8��hsq�ŅU �KyT&�^$�(�mq8E�ebp����qbR�)��	33�ߜ�?�@Ʋ���׻�R�3#Z���|�;op˶��8�q�7�{Ps<�=}��g;���"8Ùfc�L@�b�曨���CA�y�˲�X�e�]�A�A}��u8�U	'A^r���5+� �t9�#�)�ų�d��U� �,��cC}>���3DVCc�?�S���>ډ��Y�#��Z��k��I����Q��O]I��V1���/s)��"�y7pJ�[�YrٻT�%��(w%T�V��Ҋ�XJ�b��P��A{֞å/0Z�8������>,�^J��S��l|��=B��fW=�@k��C}q��X�X.����\C*��^�Gcl�=�*};P>�Dm�J��6b0Ƞ����B*�<���;f�[��ץ�YV#ԅ�{ UR*�P
���w�X_{d��o�	7]mG�m�#
#����6SW3!݈^�C����5����ξ=��i�#��a�$}������ �m�^�j��+�N6c$F�},̇V���2V\q�~�� ��V'�<,��^�(I,����w�q�ƥ��fGmܞ#F[�%�����4�Ǉ�F�s�H��U+���q�KE;�92*E4�|�+���N�K 	̂+e؞MF���"�P��k
�c���h ����\�M��O���	���Uuo�Ng,҆�Gˑ�m��s 1��M�;?�;���K��lAH]P.��}�d�m��H�!r0���7��K��{���C���R�qo$���X�
�	^E?�qxʸ	:g���;٤s��,��'�%|l�gBæ�aof(�|<2�ɝ�#�ɺ�<�Œǹ-;����ڳ�^4
߷��9K�a)�&��M|���VUtr�14�����8�O����2~��G �;��q��� ��BF��.��Ҷۈ�H��a�X���O ���o��);A[!EN�y�c�,T�'jYPYy��\T�,RV&��Z�QB�>��P�%&�B�� Y�Hj=LWR>.������ H+�� ��Tt?z���JdX�sJ�U�HP��FR�f�t��	�@���xޤ���x�ƀ'k�T���_��G��ͤ�_R��/�-��g��� �p����)�0n�T	Q���)&a���D.7S1��}N`�k�J=G�ށ1�H>Έ
�����Ţpt%n��������f6o�ۤ�A���xE�s�|ʷ���S"E��3���pgCJ�EY�E�7�ˉ�	Ji���Sy����w�[�a�e3<���e4�`&q?�$}�1�Lc~���8�Y���`��א���,y�Q��q����^r�-�<��
��'-��5�����$ �KEp*��[u��s�L��T��&�<�ؘ 6�d�0�[Eq����~��� �i�-m�o}�SMA�`H a�v�|����@�
�D��$oV�X�-����n�<�]��L��"@�����뷧�i��#�5%Ao��%d���kO�r�&7�e�k��^���D�D�cp���0���A��A�����3F�L�i�	4L+,vw��=���E��I�ˇ�X[.����r��Kp��CH�����eϡ��	˧��H�[���@���'�+�q�*�u(o�����r�[z�T9�ؒ�����
��-P�f�1�0w�_С '�H?�=�&��cQ�����𾉹��T$b S�U��M�,���ܛ)�T��bƁk�'w���fe�x�P�?���q�>1}h�צ�b_�λ8��@{:��Bz��0�^�b�2�w��4�z���,y:P.V5H�ZZA�Xq;�}�b#�=�M�#F�E��wk�nd�2Ӝ�B��[X�I<޴6��k��[z͠�y��v+��{h{ɿu$�צ�8�F���<�4y[�Jr�=l��ZS��՟8-�	�l�ǂt=���
�(�fa�`W�˜�uz�l�/������!�}[�&��� �r�Ү`�`��@{k$��1�8F�6�lB�n�<0����	�32�)�Q-g)�m�&�^4V�2	`&{���>��nȽ^�J�����Q��Ql���gI�K��_-Y��_��[�Ŵ�3E���|�g��OO��G�:BME|:�w��j?%#�|�9��2-����ĭ:�sk�ԿB�X�, �u���@fX�6'�T§ML3o3�z���H�Lx�]��?D��6������ M�����T��d�\q߇�Ɉ�n)��ij8�
��4V+���֟����2Fu�����	�NH˂,V'c��&a�TU*՗SMP�ؚ��FUf�'�����R��ȡV�Z���IfRr�#���4��6*����U�;���J�^��k���w���T}>W�%�N�J�Of YÖ_��2��r�"�m�
���a������^$��}�?�9���r�L���	jr�:����w�X�#db�<=��ηkc֗1<�B6n��W���:0B{6���W0Y?4��F���e�o(hN��~B�I7���l*���m�fZ�a�Fc�T���x�w�0�����׽=sۦ�j��퐁�6.���N�OoI�7*%���u�	�T�%
�1�Z�bR2]Ēig�T+�m5^N1{�:t��� �{w�l�̤ͧ\x�\��4-��Jh� ��{Զ�)k�s���F���<�k��D�[�������rt�H	�H#�Y{uz�X2U���2�M�|�x�$4��3�0*-y�Jd��v��i��L	^��D~T�\z���4�^�%�<���F5޿�-3�4�X�L.�xM���B�Fy��Z�������j+��0+$J�����ϵ|0������6H�iݨ�8_�6<�g�mzf����^���	@J
e�.�7�(�k{�G�F�u�,��.�C���6~^���.wP��bϋ�x	����X��3(��.��~܎�F�e����bI�J/$}�����t�<3�3��SW;3�	�����A�Z욑��g�}��E��&�`r��u����������'�����g G `��Z�Jͧ��Fo�����m����0�0
�g�����퇱�V6]�ו�.@K��|.�޻)1GL2\ab�0`Jy�=}-��3�3�!�,�ѭ9�ؓr��������Z��D�����g��t.�����T�	T	
�r(}0�����\��"�����/���F��5�����閐6��g��:���Qj�aL�Kk��%2�+X��vo��ŝm]H �䍂j�ZO�-��$1?�1R�'�ҝ�����B;U�U!X Kȩ�Wi!�G��)¥�Erb��������f�1 Ye{_���nO�nD�8\/��hw�������b�t%�:�mJuې����9��zJI�կ�W�%d娽�c�qZ�FҴ�^Ix�TZq���G �_��07u�����--�J2��lȴC$~�lI$o  R}�5�q��=�q#D��,��$9R$��7uF/��)J�`��r��\@�W�v��Q'�#~)}��p��%����G�Qh��܋�B�b.#*����	�]>�d>�!�9�\��Ԝ���>���r�H�xȱ��e��n�0�D%�$�,������c� 2�eI��#nѫ��YUI�+bF?]��H�?�Tl����ȍ�ux�D���q�LF�V��qd�&�A;z��jX�p�D=�p-hu������T�в���E�$b�Sł� �\K��x���~��f�?^��r CAG.�W���z����bג��N(��O��-zls�=�"���ZQ����RN�q���.�A��j�(N����l��Z�0nv?Ga�G��L��$���-?��k���ǌ���/����ɚ�@���p�}��˱��{��=�>;�
׬/(&(Uskb@�6&^�p��61"4`:Ma�;y��g2���JTw�q�?|�U���(����j�(BQƈH�6��d��b��\�$�}^Yn���l.��G���)v=�Ʀ�5��m�։�"#�}�UP�}q|~���U�T�+vH���������q��m��3J�҅����K���^���Ƞ���Q]R8���|��0T�"Mk�����|n��FJ�iW%3�v%?BH��fn]�k�Z��է����?])&�O(���G�QU7��;at���W��vK��{e�5�S|�_G�E���P��?IkU��[�G�-
�qe���KwHm����(�����|�x�E�ܲ���Q�Es�,��PRİ�I�zA�1
-��=h��eJ�?�H y��������Ej��I^�*v�:�A$Ro�_F�9��~׮-U3��x���W2�?θw�q��0�
\�+
3,��]�bI/d��J�jA�������p�wdk�}�D�^P^�@2�W�։�Y8q�,�-1q	�;?�v��.�����N[�wa���o�*���-�4n	�g������D@M����K�M�4t��T$[�q�y"c�-��t�UЊmjLeW��	�.�ԡ.LAo�$��&��FÖ>�w
�TE�j��,[�l ���ӱ^ gCbj��{ƫ��b����Vj4�73"��e��A[1G�d<���k�@ެ#����'�S��o��/�����%�����I�'~a�v���Ys��
�nu�Ϥ�-?dE��R�����σ���D��y��B�%�����!.�8(q,�\�*x?ڝ)����T�U��}�pq�=H�=�;��	���e���(n�B9�#R:��K��K�w���k�`X��H9ʪ(g-�{Y	���S،�r���C-�m~vóN�i^����5O��\����'�S��4�j�"`i�VY��-�U~1>6�5��u�{<p���H�AӒ?����hD�{*VgrGo��t��6�gK�2"��Jb�2a�
�w�3S�������x�'��"�����dG�����.���V'MoC諾z�r"�Ή4_�G��i�*Y0\]�[u�(ͭ	���cDl��<o��n۴���J���)��y	G��-2�A^%����5e�
�=%3<��0��G���C$����j F2��K}�C8xė�UA�qũT�H��WC�O����WmC�ު������x����}jP��<JB)l�1�8��`��s�&1��M;A{��E���dEU����cIB8�W��m�mO�ʐBf���Қq~��K��� �p���9��K>�y���pc����k�|�%L\Hv ���2a!�s
�<��L��]�"����n�,�_擄�?�x���y���U�j����aj۴�ĜT<f8��_�v�"�x����)�=
�}�0�҄&a���ΔD�[K�4���G����	g���<;	��'W=��![Uv/(��53�������t��_}�Ek}�A����m"cp6Gc�FL%L����B�]c>2���ڙ�;ϰ���pɘ^���m�bݶ�o�,|�\�/�6�E_���X,���S3�Nt�xF�h61�b��M��>�;�<M Zu�A�dZ�R�~�Y��Ǹ���灁�L	�p��17��8�q.>0�t+�kә F牣l�Ԧjz8�i�9�����CCN-��o2�����'��?�V�w��S��zUs��}�S���_�Fd��F�ݔQF���; �eogѨ~����(��"+��%\��Yf2�JD��t�!���k�h���P9Î�uS��.�k��ogi0HRw�����	�؟���3�{;�"K.�0b^օ��)���[B|�͋/
=���|V]���.+&{��2�C��=�w���H'ٍ@��dEf<%�=�N�XY��x����ƼI��z(�7�l!R0s�}��|y�5���Qi7�I%�<�T�y�x!�|���r*q��{G�_LZ�p�\O���տ~��?M��ӁD6�j�� &'��p�:u�c�飀�K� ����������n�����f����5���/XF'��	�,�r��9����,
t�{
7��;=}7�>�}��Ԧ����.�"��16 "L�R��e�M���p�"�#SO-w6f�,��4j�y��1檨!�x�ͣ]���"��'s� �|؂�`��.��ZȢ��/7�Kk��|�Z��(~���%�����3�
eIr�P�TFU ��b����@f�3����"�#�Ad�۶Np>f=��;mF/N�z�p�>�'Y7!+�V�T��w��YM+�FH[��o��)���D�R�{Z@��p�� ����w-����jp���D>���q���G���	"ov��HU���Q�) �$o1��b ^�+H<��tq�߈	4�������ǫF�Z�	�m(����=<1z�}]�[��:�����3/�f3��ޜ�so����� |�ҩ�:_`d�r���T�	6��P��rn��A�QGNv�qΦ�e��3"�?B�v�Lȥ�}I����M#��| �l�P�O�l�쇰�M�7�w�t!�rSwUie�(��σr���O�W&���R����1aW��,�(n���^dg)u�F�O0����ST+M�t��1>{Fُ�*�_7�� 5'܆/,�O�D�I��Ӏ�ؠ�U�?����O[ۋ�>p��d��M�J�K��i���0���N$��~��'�9�o��8V��rIH�����x�ÍŌ��=DD>�@3�~�!/�y�Xf��Д�lp��W�"� )j�c���^����!l���_�Z:�T�UYf���?��u�ZЏ�nN�%ك1`�h��I�y�Rn���$���a�}��al�+N�`Y�li}������w�9�qGw���W���
2�Y�t�t��T�DC�q	;	)6��H��|�=��@��64���i�|=�v��r��_ʣ6g��{1�ԥ�f����]q����ODfS�ܕ���jJ:�+���m4�l��=��u����m���Z��+��W]hzi��(c�E���C�:c3�+�Hz�Jˎ�3|���(u�"�cg��Ӗ�gY�&�p�t~�	�����5�B�\����CC0�qϻHM�����0NW�G9��l9I�� g�ᡨ���V�Q|V[o�\����6ņ���a%����]cH�Ɍ)�kH�1��8Ȧ5��g��`�_1 `�E���s&�c���ϤS�D�?���'��~��ā�U��8g{a.n!��غٝOo�!P]pK��!1�"�x�n1�[Pd*/U�3'sq5[�=��N,@�D�h�RA��dt�l;(����ˍ�'�~�R�A3�¸�h�m���T|ao)�z�q�٫�ǎ�Փq!�b`��_l��� ��<�x,1��t��x�lu�]�S�(�PuFᶼ�+��&\=���,��E�!�8۔(�$�}���O�AbY-M��QE�e���"1��\H�/��X�1���
�4��=e�Ψ���֪S*�+R	�c�ua�\K��t����i�x"VỼ��i�GW�[�ϝ4Vj�}alX���5�Y������s��f��
�I�k�bt�JZ���} c���.��F�p�q�ʕGj���#��#U����}_K,sOC�!��~���@�U��7vt����HO�l9�xL�}�:4W-�F{���eʺ��$��@9s��&Y�L�ZM{+ꕍq\��ݰ�JI����*�b�_wmV�5����.C6O��x��c".&��Ƀ��.�TB�����Ro���v7ܱ'W����T��0jo�l�q�T��M�?�K繯+���A
�Jvf�R�)!#l�E� �P��B_�N���n���}ž�Zƌo��Ā�������7J?�Ng&t���
Q�_�	'y�X�-
���k�-𹋣%A���)=�Hd@�՞.����E�7Â\�qU�Q"/�N��NH��>d�@jx�HφQ�	�2���v|�8��Tk�oD�k��9G5�	U�̖��iF��>�&cx"����l�A<���{t�8MO��F��a���t88
�n��g�H
eSN��W�������Fk6J_�GN!f������%R�P2\�=�l@ �QwL3��įE!�cG�rM�n����T �ɃDbŰ+����@��<�[���H
 2<��j(����ԛ�nH������N�0][a{鳩	Bǽ��kѻ�������ep�k�Y���f�	c�ds3�bڨX��q�V��o �m�e��K��%�y ��R)����>�P�f�<n��~o��Y��\3�DSD�T�
�ɸc��=�O�f�^~=�箫��hoF6�#��F������۱�6��9#%�Q�(r����[��%�EL��B-]y���7�����m��u�֝��N����z�+{����cNW�jԻ\�S���H?#���0/I[%"��-���ݜk|�iWF��U�hv��S1��_ؾ��u�p�r+K��E9��7�C�Q� i;w����+y��w9'��n��Z L������)��!�t�D���4V�7�R�0F����ԋR�,��R@{�[K"�\����tچѢ���i�
��x��as;*�*Q�2H�	p��#�Kժ��3�U0�Rn��k��C�W��[�dOy�Q�*o�H|��М˩W�Hp/q��E�I����һc�� Zs<�9�6P�)�c[��6Y,#؀��om*�)��L�|x��]�5�Iǟ��VV�s��rq�A����|l�]���~��������Tm�
�~�T��|Wn/y�L3�³�����(�?ִ#�u��
T�����Jn�e`�XyِJ���[sH��J�(�Q��_;�@p��S`p�n�.�\y�s������Oq[ç;Pݵ��+8�ɚ��� �!:�y��8﹉�w��G�s,W�����y����=�KA"LU�.��`5{��x�2_b��=�k����ft��#~Y�{��z�x����j�7�@���Ȃ{��l*L�tG������4u���}:�L�B0��wA(T�J�ݑ��������3L��]�#`�`ro�2���ZB k$���vv�s�q9i�5P��fXx������F�nd5;昵CaL�_B��Y@�3��|SS�MG��`�
8u��!�9SfN�p�g����-f�<L`�����e=�b�S��pqp�PZ8i8��1�� e�y���� ��g�\�V��>��1�S�J�iT�q1�Q0�`����䢘�/�[5=��Ԫ*ƯnM�rٯ���
�YP�D�	`C���b��~�� M}���@�-=0?�^'�T>�'M�%>���rK���bN�p���E�E��R��j(��W�p��@P��#�{��"p�f��Z��S�TV�u�y`0D�}�H	����Fm��[)��1��6���!����QZ�2>$Ii����*g��=3��r�������.�7Sh]�ʣ��$�Z�F��C���~�A��+����O8�f��>�E��_��[��C-v��e�������@���,)(��PN�����.$%��:�)�;��d��"6~<���<	>�2J�>]�e�7��ZePR�hR9]|��*~^������g�ل��@Ǽ� ��c+�����񁟑�McU�%Ü�_lJ� (���\�i�V�xGE��)�����U��n��E��u�8����a�^s�'��j��J�Q+>$� ~�W���=�~>�I���N����ܪ�P��8�	�)��m@e�2=tFV"�0H*sU6K8�B6����-<��8��+��In�8,2&~���-@΃e���QV����^�����Z�X"G��H��A>]�x(y
�ҫ9ʮ�^g����K��U&Y���A���4aX�L�G

 2Z�F��c������I���J��Գ/fِ�CM�����¬4�1/��ߍ�ޏ�~BT+�n��^C��9��Ռoj�4AZ���m	�]���}�AͲ��vx%#~����s�d���/|��i�ćE)ao�'�f�J��_�e��,��Au��J����Ȳ�L�"dQ0�&#��N�.߁#���B��vU�u'�?���O�s�r�j��_i�@f�@�s�:��4�Q�W�X�n'�W`ڇ"��?����9#	.��H=�GF�����f�X��d�����:���!q5��@��. Wcŵ����֋lOϵ;�N?�����6[�R�i��������hѷ�"Ƅ~T�����W��>�Lv �@I���dY����ث��g>��,1n��w�2ܕ�屘�6G����-Lٔ#E���Z�J0��uPM��7x'n>q� ��I��6֩�9�L)#���E�Le0��@G����E�yӂjJ��"�m��u�.pY��y%��U��ktxG�7
Z�r'�k����gL���{��N�?s�j[t��Y�,��㜴���V��5U$�t%����n���D�v0�Y�07@H�$�f�P��֨�0^�lL&'����]G�>B��д��Q�V���WE��􃌎j��/ �GIK�>"QE��`J�4
v��W��� 䒰qC��K,l�N� z} !�ߩ��gA����W_�rGR��Y|C�������o�#@v��D/��K QEǢ���U��d�Y�_7a)�w�Z{�~�̏�A=�����d@Lp�k���)��a��{�����E�<�=���Ni��q����ݙ_1�\���ը�PR�WB�mx�~�WU�#�(Vm���݀Xi�\&+9�?޵��f�pS��áـ����g��V8S��[��BZ�_�������6�Ѽ��%L�Yb�h���-&(k^-�X�&y��;��j�Z����@���l��]�I��p6������FD�n���b� L�V��_��/S ��Y�i� �o<�>;e��3+�1�sSY�N!�a=a�X�}���cm%4��.�m��V�g��B�K-�Q�9�"����&�Q6(���߻d�CD;1B���rz�9��=���E����b�J��ba�2�~��������R	�١#$v�<�æ7攒s%=Hh~޼G��Z7�D�/�7x#�AZ�$%�(�v����r��D��Fo�pI�r�,���!aI)��c�O̵�|	�Be�^%����op�M4{�܉���u-�k�2�M@k�_k��5�s�X�-c�	[�1�-���t�����cu��+��w��aJ��a��������k��˩��~F.m�dF@����R��y*�/i�~>�#��[JsN�F���B~$k���|E�����ƛۍ W�XK3�ҳ�uŏ^��t^�lr1i�@��iU~�Led�?�?ToYg�����r�s�5=��ev}\����a�Ug\��2 �X�Qǻ���b�`�����<�4���v8�u���^��$�s�Ɉ?W{|���1A�9�C3�ܿuS�ym=$�^�K?�~�7*
|}}��`� ad�8Ƿ�Н��^OԲ�\�a���d5[��V�U}p����������9I�а5�p?<��$$sҚ4.�x���w"_)�;؈Q��yƔ>_{g��7����;әr���aCg�Vn����o��BD�CW��i�%�SW��!�����j4 q7%��(r�x���DG�J%-���=�b5��,w��+�a�0�[��0�ٸ�/����#L���erơ^C�τW ����i��]����I|�F�D�[��#��@S9~��$������T�1�5��'gqPk��p��jı��*�F%z��n�~�x_�&�H:{�[HsNC��)��H�T��$y��(s}D�ɍQ�d.�s�b��3����);��c#��y�P ���窡�nnB�j���n#2o�FIv��xm�q��Q��@v�c�	E�f`�|x�5�����2V����U%�����L@�o!޻Dɰ�N]���Fs��y�������g�ޞ���l��z�B��H�)��	Q>ό�������kHo��ThZt�_�$�b1Z�;� #MZUJn��ŧ����Z�#��fuƛ�\6*i��ip%��i�J�/�J�?G�ܬ�g�::܆�C�<E��@����H-�&˙fޝu�ʇh!��=����3��G��Iw��C�JRˉ���>�pH�M�s�e�z�Jw�yDu`���<�DB��M�;/�a�D��d���!w�G����z
�cP�ܮ�THz�uʨ�n#W�'ĝ���Kq^��n��d�a{*3�4���B�C%*�-�M$���=�q�s�K�b�<��u�N\�xG���V��iP����k ��a�W��u3���D��:��u��P_�0��SN��;�
cpp:3٠r��Iߵ~��߮�����Q�7����k���:�ԭ��6�ڎ4;k_M���$$ Rg��ʄ�Op����6�w=X��1C�,�`=�={��T�0�R�8��Y���jX�Ƚz�%�'S��2��|�Ë��2YKP& G�"	��$��Ս��d��I��ןp|�^��+��l���@/��/�4O����;��)#k����1��՗_bH�݌fU<U�RB�r��h#��$�!G�a�����Gxc���n���s�΋Ķ+<W ���t�~�I�h
��kո� �t&�+ʜ��3)eK�o��ANZ�=�f��4�zW��jkwiu�klm�wEb�O:�UKT�Jb��QV o+�p}.�ޤ35��&�l���@	xl>�1X�}�٢Э����Q�^���6�4�6pv����d�y��X�j��!G*�6��,8{<�8���^2Q��F")pu�����	�0����ɚVO�n����!,f��c�v��^��ԛrh�C���Hi��� :����t�>�1���3 ���[gL��/���Bf\��{����k$���p���0/��k�� 4P(�byh�RA����t+zCU��r�f�}.ixn�����-l��_�ʔ0������q�Ϸ��r���،�K2b����	bd��ƕmҝ��8M�IJ�-�Js"V�GtwN؜�])'��M��r��~��d>,��cI�m��c�ٱV��,�p�o�(&A�x�$����M��m�AN�V�#�Cj8_��/�� �?�(�AnZ)��ưm�ה��*7��h�<2�b���k���G�0iN���4=g�AK�u�ũE��1��6�a��o��%���3�>O���{�����2�_�J���՛b?u�"%/>��hsڡ7��yi54�r�5W!ҡ"B�E��P�pN:f>����l��MS�74:�}�ő����^�VZ:o�f�'�KK߲��#{mP<�Y�4 \~[�+[x�]���%!c�(���J�eI�dl�yKLl��+���̚!��8��Έ��_O�<ӆ���Z �Z0�����@�o�\�[4Y/8������7=(�'a�.�vu{o"���nDZ��:�[�ê�XR�"��؜(�9�=�2<p�X:�(5�.[/Khv�m�7��پ#"��6@ eL��%3ӱ7��S*��ٷV8�~e�l�N��#�P���-ܲL5�kU���?�_S�T���bm���g�� ���$�<�� +�cg�+��f2��h��0��'�� >[��O#��N�e���
s�x��5j�I|��ꃉ��ڏs##��1�R���U~֛�~B<�`�� �w��	6����X���
�y�_^�"��ݖ�]�AfՂ%x&�7��ۋ&B^y��@�����p���qT�rI����D#E�S���K�kozy'��T����C�}�m?��ql���K$�T��ͱʓˇ��u�w�H��L���Ķ{�X���V�4�m�*�U�H#��`��d�|��z�
��*ny&�����5OO�>���ƍR�%��g;�b/ȴ�3 ����5��+wl�rs
�X�V����*t�?�xδ1N����b��1�������z�Z�ez��\�}�x��5B.)���T��i�S�.G~�M0����s���FĮ��O\�����p7��.��z���볧wf����6oJ����=L�f��P9+kS�YZI^h��-�U|�\oϱ�0�L0d�`G�"�S�)����Z��D��\d��=���%����խv���v��>A�X����*`R���ޒ������d(� =$}M��g�Kൌ���_&��@��"9���Һ܃�|��J�i�����R� �a��`Ѫ�u0r����w(&���q��fV��ʑ��ޔ��(�;��\S��?��HEKecM�4�C�"�!`:�����ڤ�O��N��wv�2�c-:C��>��q� 5�82l�O���F�l�4G� ���Oz*�Y�G��Q{/�8�%fW�%�&�  <�F$Z�wj~:��	����rޏ��'n,K�xJ��:��(��@ �I���$B��O1��j�v��o8g�_�I�����%G�r��ރ�r�J7V�f�`)T_��3����%��ZX�+WT9����Q��l�|�4p�8|����.�d�mM��.�or$
�2NH������3��}Qx�����Y1J퐝m&��N�O/��_3���,ϭ1����D��H���0!��ܲs����\��c+�b���Vf�3�e��V�B,��/���}k;����,5
�?B�8.��DE����i��v{�v�H?wdeO��?C.ޝAd�^U�P�Um�������sT�������:�i(���dљ���O*�~�� �D�b5�Z �n���X��>��i����[��y4��etK��ݐ�p@�i&@y�~�J$���_4����B϶�/D��
�W�V�+5}W�fy I�qwF~����~ϳ/I4G���z�,O�1[য���_[p��8=�ZfTf���ː`E�~�u�"m��Ԭ����!_e0m��%N��XՁ��Ŕ(�۲��&!��-���Z�H�#i\��x�0�~��<��X�S���d[��׬�`�+Ja��[�H̨+���m����eVr��M��������1��	���BP�~���Ɓ�И�"�A+��8��.�V�k� ���BX�k�ϵQ�/1^�e���'��'���Q~��C@����N�( ]�iݽl��4��+It���t)"��W�[���զ�R�8�0c������]W�y�!p�����z�ŢD�E<F�<Z��(^X���3�X�F�x���`�)������sp�9���A�oc��e��A����hd��H��SOV���ġB���WqN1���_0Z��U�ɉ{��2򒫧4�(x.�X R"�������ͪJ-�֜�T��J�����5�i
�0t���CN��_�FC �gQױ���"pbyO �?�sR��X���u�f��K��o��EE�C��T��z�Z=���Vc1�AM��NK�~��uj(�y�7j)�x�����B�D�t9,f��*B��1�|�
':n�Yb�yC2ćl`,;��6/�/
>
��h�v�MD.��qP�?x�_�Z9�)�~��F�v�4�,�EЊ���'=�װ�>��7�v��N�s�.�H��s��N}�_��<��=8>M��|���1_A6���Kw��";�Î�M�̞�yy! �b�W8A�ȡ4�^uc'�B0�j.�s�w�����j�q���F}�����E�Mq"��M����9��\��`�N��E7��� Z��%�++/�# ���@��+��K3���tMeZ�Y�����|L[-&��^���Q�ʐ�*�Q����s��!�d_*@�i���c�zR�Њ�}"�E�\9Z&?m����W
S�Ԧ5]��co {l&�SnZ�a >�,��+��	?����(��ag���B��j���)0����޳b����Y��k<�a����+A�Շ�_�2Q3�찔I������B��]��}�.�;ؐ�љ�@�a�E'��N/46��f��t���ujH�\�T�˜^"�~��&i� g0� �޿W�����p�����O���{�oQ����%�����a��.|���pq֞�G+�&_i�Y��d�?a���H]d�#�Y\<ϵ�� {^vz*�5���M���S�?��T����l�InU!P̏W�r��$ŕ��z%W�o2�p���
��L:�1�? �K�$n���M��	�Z�"�+FD�y�",�靷�54Z��'�'nd��Ⱦ��A%Z1�K{�|v�h���my�M�����Z��UȻ�r�H�Lݔ�,C���?>9�,��?�W� ߹fr�����Z�P`<R��u��M@�RY>^d��h�_���<{�]w�~Q7Ѣ"�k��fj����b}�E�J�zFz�e��zV<DYp
��t��uO XFB.�#�?әXyᘛ�Uy��2 �k MZ��D�J�$.O��Z5�(,�7][���\�|�;>8�����n�83�+{>}�\"�G��ʯ�2X)m��Xf�-Q�ԯ?��~�����Ih<�3�N�P��A[�����it��P�׎����_�m�9�X�tL��0 h��+�'�;�<lރW��K�����@[�,����K��⊻�/�	��I9�P�>d�´.{P[�<Qx��^�G�@"�&�a�4�m�3N����a}N~8Y���t.��(�g��Ә���~Mr��))e�j1%�<��N�� �o����Ͷ4l H�+���2wΎ����-��tZQ�F`�3� ���׺a�!�����2���m����vbY�y"�k���|{�De�<������V6�C>�� N�4�?G�8]L3�dm��Ũr���tv	}���0��ȼ�M�vi�?�����*���Е�l�OȀ��g=g`�����ւ���*c�ma_{>��J�JT_����~J��W\�{D�y�P�,A#e��.�JO��K��@�xKB�ʻ@����}�W\HUʂ�LDLpk<ةcv��a�_+[��{��%�q�ƙ+^�x<�e������]���FN�qf��a��P���P 6�d�z�����"�������{y忷����$r���E�G 55��\ ��[�;�������������v�`�Y�Kފ%p͖�}�ɮ���Q(L�D�ؘ���Ʃ�}��My��eIʚzH��R�
��"�I�Ю��_@��v��ߴX.�$���F��]]���rm
��O.U��w��*��B$���Q�GPC�8�N��xT�}g�[۽�U�rw55d�5B�a
5(�N �v�k}�^�D8�q��')"�{�N�Rъ>	��f�S'``z���;�g�"���5�S�4b���� ��F�"�i������������}J���1xj9�����<񑳎p��o`���Ӹ�X.CVTU�%����=v���8���E�6�ΰ��b��~���?����Ʒ�ryN�nݻ�]l�[>L!�z�3��-/y�9����;Zww�on�#e�����-g��v"����LTġJ(���a$ �����׃���]̟�_��g�7��e��$RN�`�v��?eB���8w�k4C�GG�!}�$��yy��_��`u��1�9b�a|��U��rg1C�9� (�;ˆ��J���Rc9ETO!t%�����W��d��NE��-S�#��P��E!�{�vO�n��R��W6�`E��_��TXRS���>e���⡤Ki{4+��	d�1U�a�w,�!�(A��_w�GKd;� .J��.��	m��G<�f�_�ȱ5�<��(g���u2�FZِ��!a���ފ��߅����PJN-̼���*S#R�w�j�u� �%!溹��B�;�f֩ՓMR���a[Lî�̔y0�������ا��D����2�:��K-����͆%�0�Si`B~>�w�OV_�_�sSPh�"�#�$%�>�_M�X�<D�@��'*��ہb�H�|s�����Ʉs��/�*���F�!��.)���|��k�5\@L�#���� �l�Ϟ�і�1��.�S��9%@��P���r�;��f%����g�s.c��Cgg����O�A�4N����2.�Jר�����"�M.�i�
���i� �t,2��Q���`��N� XU؏R�Y�E_T{��ãG���_ɦ2�n@.�LV�3�~�i��:�x��ݨ��Ɵ@���X�F��&�j�\�e��V���k�|W�<O�,���9�ߓ���i�fP� ����)�Y�+���>U�L.�[�<�i0�%���ʄ�|c.�#@&�=ӟ}w����7x5h�s�RA �󎔶���)�.�,���i�5`�s�k)� ���n��.��CdIa�7�X\\j4�-
b$nkmA3��W'�|���������Z���Ӭ��VZ^��F�4p�b�����<q��I;�+���;~ПKD�����~���8R����Y����ޅf>!�+�J8���&�h��� G�}6}�xa�GwO������6�N��%���/�����~�o|�r
�4�H���$��7���yK;2d�NN�W�Yr�/]�I��3��
qO���k-��W�.��o�pa��t��e���e�t�T�愀0Hlޡ���G��s�� �ń˨�\��'�KiD��X 4K X���;��
Ia���IP�E ]��˂���TP ��3�	�\��a0���Հ-�m���C�X�s# 6}��p*~�+rTM)����/æ-�R��M���H���L��������!��%�y�y�M@��s��������k�������$��m�r�D؇��C8�c��Ő5��,����.��b�3\���7�v����+��A$Y�IT� �p��}�k��^4&j�و�K��-^J����Ğ��������'z�0 ��Y��3��Ww�V���&�BM.h+X���Yε����X*�4���D�K�%����Ő�c�p����4��p$�ǈ��YR�������W0�pJ*{�c�G��k��9�z�i��+��n�u�y�A�m�	��
�-�bХ����;N���0�ħ�4�4Y�$�7�E]<<�c\��Ҭ�������uY^N2��W�:\ЕmSWC-�Z��,ǽ( �fQZ-9�:�a�a����v�e���I�vD��7��t�v{S��<�Ρb��7ge�ϊ�Jt�I>DeS�2Ͳ�~�;QsӁG\����g/�3����I OL��,��ɟ��	�Xb��t�!��b \▯��$b%:9�3)�y�|��)��5�8?6��jr������q����e}����M����-8���Ć���Z�$����<�ō�l 囎�������h-O���$����la`�=���B�|�p��{M\�S�/޴���y�s�W�l�RGsy������/�z�����&�G��`x�:j�u�������up0�:H\�Kf��$",l��K�����B�� ��EKJ6O&'��CE�ض����.��Jy��wIdZ��̅�R��I�'v8%�J�W���� �Zw����O26��<Myf�f}1̳dZw��)E_0�A]�>��e����c�RH�N_�Bz�Ƿ�� N'�_u�1܎Wt��uv���F�W�||�n�G��0X��os�hQ�W���y�ae���6blY�X�Ju�ґn���Ҝ��������H�ª�S�� L���KG��`.i�-�κk�W�@�� &��ջ(���8�kD9ɶ�<p�?�>°����U!jf��|�S�H�@��_4���E���@��2 )���N���A󀍷> 
7����-_w�@�� =Gة�h1F�"e��;E�� �e%�r�l��e/��J�:F1�@��UKj�n̾�)��sI�����/G��h��,C��ц��K
0�q�e�P�"(-��i'`�y�6�H;�%�U�X�k3/5��	Q$�3��n� xK�H�ؐ@�6g�������ZE��"_7X���fOX���������L��b9��˘gyJ"�O' ��R������
/*����;�� �Wn�ܒwvL"�ĸc�k�LoE����ݎz�z��q���NuV��^��sVK��h:�k M~h�lMJ���^�?h��
w��s^ R��D�H�d=�x�0u�+�3�����Ą��Q��Rּ�os�/Ϳ��؄����fX|}=���-���y�����R�3k�
t�vl6%��I6��lj�~gDq@���
�yLYZ���aĽ����/���)Q� ��Kp�������3`
�㾎��
p��؁�OP
5�	GޘŨ��}�%��p���]���1v�u�T�d'��ɓ��	#v�#Y�6z�l�tۂ3���D�L"�����|t&��9��r�ey�V��7H�C�*ޚ��;H��㵁
�(�3m�<N�t�^��	N�+���eȁ\�R ��o�A�����!yl�^eJ]�;Qe��Z-�2؆~��'nv��z^�Ȋ�k�f�:�#X
��~GG!H?��e���(�f��C-��y_1��K"I�q]����8ѬR[�z�2I����?D��\�%�OIm�/-}�Hzo�ӉG �N�Ni�&dh�7i΄?r�w����)`�*G�ށ�?�x�ec�������&�Ȯy�̝}��񷇏�2c��������6�i�sH���r��KZ��|'�>�)��sO@���*Fa�h��ݰa���d�K�;J��]��&]c���%{�I�8!��p�o���Y��P`.��p@��J.m��ޅ��W�B^��*;��Tx�pq
�v���ʶ��}ќ�	���2"�g��W�x�<�Wx�s�dh��^���K�35�gg��\ۄ!Ŝ���Z�ZnO"�>�цE�/W�89L15̩���<x�7���f{/}�0M��+��ަs��~�T��f��	L���p�%=��WZ��W 1+��h��;X��g8@���	�^�jV0�{�^�yb³�w��D���$>[+>��?cxP��R�`���{V ����(��m���+��;΃N4ޖ8h�UX�f�<ɟ���Ŕ�[g��'�:�R�@��k�[��@��z��O�}{к�rV�$�2�U������K���Q!�I��9�.����������Ztp��V�&Pp��w;��j��o�LBĮ~p󮜖"6�N���.��ըmG�ݟ`F`ԛe���q├.no|�6&3�f�}@"V�V���/Ezm��Yye�0��t����8�%I����q�(A�X#·M�4��{p�� u侹'q�J�p�zV-E+�����A�N��`k}ƃ�{����u4*�3�Jc��zq��@����!�(���]w��`�������5X5~XIm��18%'�	7��r�[�k!�u�N���<{��mFО�9`0L��|[����F����I\�k�P�K�S��j,p4D���.hVң����ˑp�eB.�ŀ$"�0��{����N�����:-�J��Af����3�N�8S)��@���S�ߵ��C�Ao]_,�φ|Jॷ�{;Ǩ��YL�[[��2�x1��� �3�`�j��K?m�o8p�{�*=��?�2�R�m֝ d��s��KU�F��mJU/_I&��5�U�5��qm&���*0����ZX�x8=������ǘ�Vӟ����B����B��H)������6������ٯ4,0~���sY�����*d0ڡNJ-_46t'$5�^s�`��KurI抟?T	g��ri[]�,�s)S�w{�؀��x���s�Ⱦ��i�pf��������p���bZe"��P�_#&\bn�i@.�]����ာ���@Q�����Kީ��%��H�l��&�G�u���>�OV���V�nJ�
W�����򰏌�I�$~a�hdf}�a�:�Х�6�z��S)��${X_S� "'(x d�~