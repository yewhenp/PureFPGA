��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ� �t;l7�U��ಬRXܸ����ڮ�[�d6;�y1cb��B��G��d������|L�����4��MK��:��x�j8��'��.ϻG4��-��iFY����;ո̈́����b&0d=D���ޒ�%z \�J������P��#%j��E�I�f-����9�<�J��Cث����J�Y�6̦����2ڗ��7��w
�_r�M���|93�������P{��M%G��\?��$m�y� I����#L�̤"jX�_�n�ޗ���!v>�|����Wg�P��7�'��4Ew9}|�v́�cI7P�7�����%�y*~��k|/�/)�y@M˩�!��ˊ������6�2��׾���Gn�I���G`Y\kV��3,<9�$΅��[�Ui��LIQ����? �in3Y�����^�U�3�'S��������p��������Q#����͑�TT���D.����{��[l��V�s�䨕=��R������/�焄�] �)���
N��,������~lg�lh�G]�)]4)�m�*��(N�L:ؙ5Lj�� l�Li�bF��7�����*l0p�ÿD߷���Z(������w��@=̻j;s�*$.�r��m9�������h���:���~�њ�	ZE.�ϐa[ѣ��i��(��$�lľ
:��C�g���3�9�����Id֪݉�[]�b�d��S�X��Τ�67y.���)Jn�j��9R $\)�2�Ο���)��n�r��xu��qoAP}h�5�6���?�	��w�z
�ԫ�q�{�ԙK���f�� �xnMS�hy�4˽�� �e���re��&�I$���X\>a��\N~*;ي�8����sɐ$
�Q%S���R)p�3z4�/��W������^_��.��OQ{������aRS�0������0�N� �E�TA�@�,g���?[th܆�/I�{	���.�A�������	io���r(I`64���d�^O�Ǟ�r�.��+�H2z@b��!&8%��a��-ղ�!�
�H��JF���b3=�ⴒӶ��䠬�Y���\?N��<%��&k^-'��v����R�	�T`-S�`����ν"���#a�6a���z�*�py�b[Uf�$�W m?�#�DD�|t�ۑ�6���P���jN�����jv�>�싢���
�G�^0��t>����T���}.��]t�F��L�.Ph����bI�o#��ꧥ���R"���G:���6p�$�ng1�wj��q\���o����cT�zc�cv�r�;�����k��B4!\�g}M�
j���r����@V�59�T�5�Ǐ���v)'ö
�׷��)�*�6�6L"��͹����.�Mg��h3�]䫉�CV� ��6D�t�'������z3�FG!@��i�S�C���͹7C>���!ʌ��"'`��xߕE.v��@�*�6��uw����`��(�/ER�8�Yt�k~Y=Au.`��F�h���DcMg��>�o�	Hde�6�ER�C�Ѹ��{�=��B��B�J	7&
�f��KV����d���&������A妨ΟH��P%=$�f�/�����	he����\���*)�9��HiX�;���/���|-F�!'f�!�L���z��7��Hk�Jf��p*h`���Sg�DH��A��O�UiI�$����,��{c��n�S����1�f��X�!�#��k��N� A�
g2�o����ף�s-cͅ˰���s�>~���K鐐�-xB��{C�F���K�MS
_��ʯPt�Wz����o��m����s89g͐�B�u U��8��C%������� ���wtC��9`�'��M�FJ�m�ؼ&<S�����72j^
����z�p��s�U�1����H_�L(�����u�^��4�Ό]e�гD�6Rtnt����2��Yu}1Â)G@���]m�n)��ܬ5g�H�-��	�}-��w����*/����t�b�,|��f�W�v��{��}C�Ό�x<���7�f�N���Ї�NO�Y�R_$��	o�������i��'��,����?^ic���w7�@�}ѯ��5��{�pВ�u��đK��xd�T�$��*�%K�e��?�PK���$&��-��L�G��v������,���j��� K�����q���-��S��42Ĉ��F��s�mW�of_��N�MB�y��_�~2�0��4pK{H��0�;Q�n9�]OG�8�y����Urk�� �G�+mWx�4�O�r=��g�h#WX�$ݓdrΧ|�O@h�T��IG�ɮ�C+�ӿ������_Z5��	���}������$Zx1��A�l"�̅|1I�AS$��Y��$�|6�*	P)��l���@D���ͧ�"�� ���H�n_�w����ӵ|#����e,�1��R4��<�:�)������nK9�S��h`��/R���jU��=�=��Q�N��+%�����_����$�@g�v�p�ӎ��Rc�A�
�E7؜�sF�^h��ɒ j�@7"�U�G�\�!��06�i��=0���3�3g��俜Uf��T��K;r�9�n���p^�DTv�	�# ՠH���K.��c�C�#�aZU�q��eZ�w�d����`?6�l�[_S,+nrMsZ�k��l����o+t�E�
�<�9�@�����ơ��8�/�bﯓD3i�AW�W'���R�q�ϡ�M#6�b��	���?�I��T�m��=�81ϕ�MS��2�*%��o�53�n`%Y-�5����}�8�0.��3�)I���l�n�����E�zRoOQ6ݪ��^w�j'B�S��ޘ�υ��Uk���q�Ik��R�K9K�W�ݚu��nf'V�QJ��|����_JE�ɜ^f��;�B���P���jP�c7��*�Nmx% �f���1��,ePr�-�`��).�D��J��v$��n����~�D"�(Y������}$�lz`�����m���y\@ē�mk�J�+����W�v,�(�x�����f?�Ck����?0��Yme�4��=b�l����ؼ���q��_�Ǆ�թS�}�Q	� \�%����Go��h_�^��~�_�|1${���\��w���Q��0��� H���Ղ�ȿbA�nyM�r�%����wI�7�[P~XǯJ�]���������R��a���ҋz.<Ys��*Y���_����]�q��d�E��b�8��Ǌ+��8U�� ]�ۢ��̥~*U���yqe�R'x/����ն/"s;*�9pj���h*~�`p��q�P��c7�]��#?���L��x BW���&��1�R�5(~-�x�dc7J8� Bx��������4j�!���R�c/q_jb��H	q�E�����{��k�N�L��̴���6�G>Io����I_Z�.38 N|�s5�q��ᴿϾUOKu��)���\��k��g	[�S�_ $�(��c��'�Y�Q��ªeN�K@G�͠��Ek3k��6񢹋�K��8i�dZ�q3��qE�3�����8���;��}$)��3�i����A��9p,�@�-�?a`<y������a�o�N�X�'g��.�@��ڻ��R�@��#��w<I&RP�GW�D����2R�x�Y� ^��9��|���+�W �!��T~ z�!�X��+�����4�u�'�R�:��C4�#y(��#��Y�R����8��g�H�Mu�����I1W��c������p�f9�0��y��d�8�yn��h�[�3���J�_�� .8�t$�G b��0�-݈�ws��x�o�uz�y���͡$��Ϧ~�e$q��s�,;�:%��%����cT�Ng]�C��b��C<��M�j�Jk'{�Z����@�Cʀ��9>.��@� �;���5v�������k�[��-ؑ��{�[�<FV��T��� w�XMߴ���dGQu=yB�V�6�����՞�M�� !48،�]�W���4�6�{U�N�b��a٬��ł֑�U.LAQ�<��jѤ����-�g�9'��[�� �$��b���41V}�=K7�t��c����-�DN~�$6��'b�-�����w,�=�~˓��W�� ��~#*����B��ƗL;<0�\K�IITS����˞�|'2QKIUV�X�'q��2�6��m(���T�hP��[�u�LP��o׷xUF]��TtLn���Ns���ט��i�Y�e����s�5x�G��Y�4i��<�l��YabWar՟��c*{&@g��j�3EB��8�2]Q{{���i�j(<Y���p�GG�	���,�S�]� �Ý�[uG3�-i���I��~�2Ռp<y�"���s����]�{��C������GǋE�q�s������Rԉ�a�8�P�直'�=�o��y��p0pqSa����E���'i��D�#@?���ߑ���/P3D�۷p��*�&��N�ؙv*���*o��/5�"m��p�vu~��?<�� E��AG-b���ϿA�^��n��`���	�:��^K|���Uq�>v.@�R���YEYj3�����uu�=!�ث.,���;���=2��� ֕�6�-�k ��8`1�C/��]���� c��1rk�.{Jz��\�j3F���;i"�����ҙk&���#��k�fS�J�g�Ϯ�(�n�$�F���!��rEE�>p<��'2��d�>����_L�㚨�q�.��u ]\F�GLd�n6��Ar�GwV;J���@S�ٓ��ߏ�*������.x�+�D\�B���ж�:[��yd	@9S#Q\��a�!���L����|�%
�	M���9�
s�w&��[���Wl�C%q�&�4��54p@��|ې����;��CF�7ilD/7���������i��x�(o(��|�Ո������4#��Fvd��`2/��8 @��1%����-GW��V�v|'FN�t�����ɝ���+���Kp%��P7-��SF�ɣ�J =�޵c��8w[.:G�6�NK<W�U�jºp��qP��əs��Cg�,{�t,��Ø�%U�}��/Q���B:�l(���h��CGN�,�p���OQÄٺO�@�N�U��xB�arY���Q�Ŧ*�r	J�`���.�c�h���{��K��D������7F�&-uz�x&�K��&+rp|�	}��jR�`�{��֏r�l�ə��.opG��Iy7�)�.�(���p�n�gJ�]&�,d[��p�.�/�

�s��*�P_ċ��?.��� 7i��f�>��M��֚�d^�K�_+)�#�A�T�������l��ZZ���ه�#�3;t-�K ��P�g�n9WX�m��/G3���"ާ��SR�ԯv���b�FbQ��v;̀m�2m��L��U}�/��|r,!ةZ��|��2c�a{sg\��l��!�̖g��bW���ʫ����يX\ V��ً��ҢݍCe�7�R�����Γ�ۡ��Mm��� �T��]�������;�c�� r����\I2UY�:_
ͩ�h���U�W�� 3S�� R���[�V��~sqǧ�}b2e=�v��l5���=���N�Q�A\7�9�����8J��A�Gl�o���苢�,�4�4.9*���s토�Ed{���}&)����<uXj�<d�Ys��K�CL���+v�sJ��܇���pZ^��ttZF`���੃�a_��Ơ��uϊ��*�� ��%Lm*��=X�� ռ�?�?�l3g�Ґ0<u.� `�r�V�V*�c�ƬB	X%b̷����XAi�~	�m����Z�|���I����j\<9�Oe����\:��������X[>�P�-rD/Vݥ|Q)l�	8����z#�����g�aI��b(��rս#{�C�K���!2�1}�؎j�In	��]s�N���XՋё�b������`�5�ɾ{5���;5�Qq9QLJdaӟ�Q|b�"���ՔU�Ҩ���-�S��Bä�c�R˚�;Q���B��ѺT����;^�MҸ���_1�1�^
��ycr�Lȏw%p�a 2��[�\�:��|�S�Τ��95M��1��*Ypf�YY�׭4���T@l�����s�1j�0U�I"O%Y�H���/.���"���֧�i� U�#��$�#6aB�6^.gy����� � �N��%S��38;�l��O5Qq�b;�:���)X�J@k��~���.s���
/6�A��X�����f�(��H�tݠo˸N�&b�д�v#���8�j|j�'�M��\^.�^�sok�?/���:5+=;��<'uԐ�Rp�A�1XF�.I
X��@��l.X�C�j%����6�;�D,�)Ι7�\��q�KC�E�ٴ�`�ſ������ ZH݄�R�<�����8�S4'GS�ߒauHVȯ�]ç�x~P�p&fZ2]�[��X��O��M�O��)�6��B]��P۟�]N���svR�o�/XM0��F�*�<|�Y?�P�/�׽�쟝���@���(����;*\'}	.� �`�$�]8����9�(���6Cq�X�jJ�B\���l� ]��P��	�b��7�d� 	.e��^���%y��GR���Z���K��;���2#ޭ�+6���!����ȇ]�S�vP���N����?��N�Sߨ>�h�;2Pq���p�6�����,�v]�M��6�)���\n��0�9���W�Pے0{#�$-,c0(G몤���#��P>*5�8f�7��~tR\��+ܩ�V3,K��{��3o���Alw�b���:揂�L��a�ZT��g��Q�2�05���y��+����wjƊ��$C1�u�05X������wZ)��A!����ž�<�!ta��'+�Ǝ��Ps�~��*���8>/P��L���$�8<��n����ۗ	aTA=�]�U<r_ٳ{������{��-J�je���S�h�7�m��uf� �:]RU�?٧G.��֡ �U�D+�h�LQ���S�GME%���$��Bk�=�̒�!�%�>k����B��{z�t9gd�ή��R�&�4)��q��h¥����>��|t0:~n	��p�b��ɾ���<>[��k���p[�>u|�lNw�y�ӵ�_���͸μX�ɧf=]���Oب휚� ����K�yf���`N�6^j˸�6v�NO� vȼ�6 D�-rtw�v�i{T>O� �#��
@����]H���������a��r컀�ltF=�׻���B�T���C�X9||h�>�-��c/�e�>���+�O����KE8�Ք��XD��O�?R�Ѥm�8�I�&��X�{"#R
�b$;��� }�@S��^V	�I�l�K�u�C��c_Y�@�	OL2��BjW\l�e���(���尀�[xXQ�	�����mV��)�<M�$I �a&�n�)��_^}�_^���ABz����A�E|�P|��nw�!h��C�u�F����ז���~r���C	U��e�y��<'(��n���ql{iC����o�������iSV��ͨH�zr��B#4���E8։o�+�>s��Ę�;�ί!�@��B1W�r�����|P�P������ӇX��x�ݍ���a~��@6Hf誖�<�x ;�g8�D\��^�͑	��[��&*�m�7>���R���fe�����py�-|��K��/q)�����Ɏ��i�o}�8E�Q��Q�;]���We)`z:lX��\��i`R�"^��*�0�$��[�E�����8K�u�j�03�UW/�2?d��]gfMIT����%o]���$	聜��;�8���oj4�8�9-~���l�Zߚ��)�}���4&�ˍ3χ�!�o.$c�|g$��h]d��t�"kHc,cÐR����+T�0 �����4��C��}:2%>�
����Ti�(��!�:�7<,��Q��7Tչ0;���?��[T���lX.g(1� R����	PP�_}qU��&� ̓	4��5}ږ��myDH�����V2�rU(|�:^ߌ�a��8T�1���T/��\����-R�˩����Ő�O����aSG��((A2��nG�ױE����u�MfYN�g)�<���y����6ZJ�Q�#g�0@ ��3T݌�)|6e*4䷨T�k��S�0�&��}�Ձ��,��#*?��������;$ȼ�08��ߥ��C�������4�Q�o�CO��h�H��4�s�2��a�m##[`����'�O��1��N��@���t�
���H�� |ܐ�S��F�Zx"��}^����?����bS����\�K'd�An���,��� �s|./�����"���p^��'+��Q�ӶfR���j:)s.������(ճl�jU@R��=�Y
YuI����0.k9�ǟ�&.I|cYa�&�o�U�d�z�_K���6$�d3T$�|�'{�-�	�MB�i�ςQ|���f��@�U�m45�q��#̼[W0s��)�,�\��Q֦q�*$�j Շhpz�L-6*ę4(政ͭW�������O��B�s�3t=r|��~����N27�/hA�VJ����#�*!���=��]қӈs��:�e�w����e�ϻ49+�/������������7�����Ek-�JE?�,�����ŧ�t��bP@3v��c����6l���t�'����u!���0cF��^�`mA$Q�o��%��z$��v�;j6_0�E��.��Ùd;7������2}��\�$SB��Uy'�������Im��o�&v8��v���!%��U�%������˿�
Y�n�O�0��C��|�����H��Q�����<����D�����0o�8z��G�8:�O���e��尯�>x��V�ܪ�Nt02��鸺���5*Z5Ûa�]؍��
��2ㄋ��:���˟M�a	�� �JU��d�V��z]
n^���s����q^%9Y2bv�sj�ZbE.��TF�(I�6J�/J�#V�an��ӳ�����ooo��D�E�@^�������,	�ˑ�Zk���pR,�Q��Bâ!�S
�ް���>�Ȑ�h=,ls׏�U�!�Z?�<_%��^r���Ӄ�ظ�y^�'��\V�G������Q��������˶^H���[����]���lh��k1Y���f��z�\h~��@�Bwт�^+� ;��O�
�t��L(� y�|/�h�*��5R��k�RJ�����*{��k�K&�� &_8䱸N�2s5n�Y���Z5�L�(Gۭ4���������ѯ��;�C�E`r~��6��۹�ړ@J��ӁOL�(7��CP�z�o�1S!! �ʫ{���8���D��g��ik+e����]ȴ�g��M.�?�����[<>�3�6��<���cN=�ߎ<&�78������m|�yL��>a
m��AĎ+�t���Pi⥇l�i�;(��!�qe�jN���f��V$�F��hN�&�L�:�sa%��������3£DT
��~�vn��!���ڿ��-H<}Ou�~�囲�7a^S�#�8.���\�i�;��~��^a����ȣ%^�r��C�Yv���/#PM�MȐ���
�NZ���;��ts���]�E�w
���AD�v��=j��2�&8L�D����,%��3��џAyB�3�QՓ�jljKn�C�����뭢�F���(GF=l��n�87|��L�+�=v'�.h�����7�m�,^�����2Ϙ��~}��Ĭ�T6�!T(h#�C�+d,��n�}	ϕTW��Ҥ���ξ��ȳ3xf��:��<��Dj����ط�~�����{wf��53�¾�D+�#�{2���(�
��\m8���E%V��K����+Yl�FJ�N7��U�T��!l��b�>�l������w��_����H�,Pv���8kN+�'�����������U�h�h@�~pXB�}����iO7�9��5y��q�Y�	iq�m
9�������c�{��7�fP0#/[KєU��4Xl�xg�8��A�{��0A�N(���tD��}@]�+:��piq����yeY�8O�D2�H�(Ny=Z���ɴw���b]�/滋X��-�Eg*4�j������{�	X�&�w��yL�aj�����S<l��N�N��{t���Hd�uf�B\R�L�kN�)ĮI�B�)�o�����9߫�;��!��F0V��~{��Q^�B�P�w7kMEk�K��~%�� �ƷA�8�٣���g��Tk^���y�Bt�/	
�D��q}q��e)@��z2*�;5�Cb"�ǂ,\�t�L��EH��z����^���4�Ӊ���6V�\({U<=f_�ƾ$N�S�&S�g�Sai'�Z'Hy��W�����S��d�;��wdCN�6�q
�j� �/c����Wz>p�	r���`�M��0D��� �~5q�B�A�3����(�s���W�?��O!�񔃗��'� 9���tܭ����{�?[�J݆
�a�\�y�|�&�k���/��v��_�A��'%��z1͈��:���S�h���S���{ua?#��l�#uᢨ�GJ�̋vb�#� l����vJ*�orѧO�P��F�s֌���+���|4'�,Ok���o����`��乕�W -�8HC�L����dLء��Ʊ|��QF5�w��-�o������mlOb�+�D��U^���WG��}�Sۀ!eQ҉%A�>����DͣL��U��qxrB?OҐ~D�oߥ,�z�Z1:��1�ʭ��e|�c���	����R~��k��e՛X�E��أ�7)=Yk�&\�1 ����p�MB��]�-E�i@VL�r�)�Tq��X`E��?LN6�5(�B3P�[Ki�鸦��y��T�t֕���ʂ����`���9����&���,$�H����������>
���D1NP����z+��m:΀{�#K2j�o��_Ve#1�W��(�����9Ę�t������3���D�x�0\`%�|�H8}]��������F�25)��FbU'�=m�BRY�&Z�g����U|�nB�fzC`��=�F~���~�O�|�!8:K4j���*ڤb�ZH7���/��lT��Q)EjC���_`i8@�@3:�w�[7h̟by�0��9-�O�m�F���Lû�o��U:�Jä��.H�!��EU/�F�Ŕ�)?�)�]�U���M�iT�3�(Ϋ܈�o��<eh���0�,P�נ��C��tAY�߇I���6m����^��;- �,�P�r�����������۴{ݠS3�ۡHR�3�5����a�N6����t���zܑ��Hr@��Q�PΉ}��XS)�T�a���'��+�% �F$�z���\�fa���P�eG9;W4z]��X>��O衳*�z�b���5� $�V���?ީ��S�l��~@`�ʯN3��1"�w����[/��M�AmK#�p! �w�XG�9��!-�A���$��%�hˋ�WS������ȐysW�;�8�z�]��|��2%v��B]{�H����qp���nt2X�bW	��%���Te׹��CdP�̵
N��b�!��/�挾�2'�=>(ޯ�\�{^��+j��g �G�:��������`E��憲I*)%�4!�#⌶��Z�I6�R��VWغ���Ez}�}�v���TdǮ�k<��2��f���Io_���<��Y�BJLƆ�O4��qw�(���g�E�X�y\+(�?������e��[� :7O��ȵ�&VQ�1*8n+:T��9�}L�߀͸�����(��������@S����G���8����x���9�Eld _�I<Q���ޯM 0���aآ�������R�8����bB�5��Ŏ�d�P���\|����1FY���gW�"�Zp�~�u�#o^	+�rǾ]���o2�_R�̤+�&�L�;�kZ�T��gt�Q=k�*9!Bs�u�R����W��/<5U5��(�;��HӒ������s�?Kz�@<�(A���[5�\T׍a����>)Ek�����{��$lӚ(���G?mn,0�|a��^����4_ڟ=��l���knU&.�-0 K2I?���4_��������G_�&�o�Q u�Y}�l��Nޟ�7[��7q˵��P�&lJ�����1m�Sz�|dQ���Fv��p��D����
��!�^%s[We&�w��;��O��7C/�j���;����߾�ݥ��>�7e6O?�
��ؔ�Ն��?f�a
�]'gU���
�}����[����|~�k�Ֆ��iU֟[���H��9ce4�s����ת�R��1�4��4q�0-�n�d�bso}�Ɉ]�빭J�Ƨ�l��P�{ZU�[2[W�������Ɇ��Ͳԩ�ur��؁Ζ�x�4��N�I?&G���X俬��,,�+E0J�D�nÚt���&~jU0�b%�\�[�lN'c(������ô��І���s�>W;R�|͋���S�gj�OS�$���p��=d����B���  5|K��G����Ȯu&��dbۯ�Y�wλ���v{��'�-������D-��L.=�]�_{�.�|�iSUpYI��K�Z�vh�\���s���gC�܋��s���4���B��?M4>�g���8`E�����*��"��l)g�
mM�t�-<)P~Ri������ƛM~G3�E��o�,}��	G�̯��������~�=��J���a�>�	W�Dѝ *����gc9��E:M��d��{~�K�t0����RX/|'S:���+%�%�۹3�����D���������Ù�h{x�};�~&̵�Cd{���h�-�=��(Ϣj�n0D�w �W��m}��u1 {֦�!Ʉ���t�=��8��sSm~��bׄ�չBFێ�ٴ��{2f �U$�����*-CQ�
��x��\ɬȽd  3��g�ń]R��`�˘BT�Ԑ7��Kf4:81��H$����r��3�LU��[�ZI����:0sMI6^0�Zp%��y��}�nyb���`�O��ᘈ=.�9H�Vga�X�~!Z�e]f����!-��NQϪr��7)��t5}�ā��)`�z��VQ�-�=E���Se�m����\�B�(	7�d�s��;�0��G�+��!���q����@�!��T��o�A�C5z#���*���8E�'�p�|���ר���hi���ş]y�{(gO�}j��q�
zteA�w�<�ՠ�qa|��� ��R~}x���1q�c8{ڡ�
�kؾ줯,~n�}
�فz[�m��#ggI�����E��ؾ���
�"��Y�y`7:�~o�me;���tV5�L�F��WT �����&��vj%S?�܅�^��� ���wC��ZrT$m�ӮS�=xW�i(���s�O�!���:avha�v��`�ڬ�O�):��4�t��mt�j#V�ucU5;&����,V<�2��|����{@�x�b.eO��E���R�_�I�����H6�Yt� \����'�ɻ��EL���\�}�<4��wB|eݐ�����m�A��%�B�w媉�����}S/��?��c�?�?��v�B��Knb�1(n�5t�����9�W!�QV�'x��:�>Iw�CZ���is�~���7��h�Ю�D9�@6��a�
=�/�UyƤM,v'+�U��[���ſ=���������;s[��^���4�g@�!�=4_�����ȪÎ���sh��G��l�p�߬�������A�HҏR���=5��߶p�_ͳ��w0�
�ˊ��6�e��(��;��yfx�����(��)�^�����fֽa��d��=�3��'��nʷ&���'���ݧ,1ћ��}�^�.t�b�n�7�O����no��*�G�=�\;t���'m����2�.t���4�F���%��a)k���q��
���p��CyA�hJ�c�S�n�
pK�LrgO�p+��|�IJ���tC�g���uZ���(���>��&�"�xK��L�# �f6��O�*�1�#<�}C���Z}�1�<(��7�\������Ӧ�Vw�?º�}&:�(,�n�T)�.-����g�ޓ�ln%�.~��)��b��.5T���kRs�_db�5A��{�`O��8nɻ�}��P�3®ڂ-w�v�7�\��j�\��DIZ�$�>x�m��鑼�K��z=�el��*/MF7�Yet��vzB�ȥVw�.�D2RC'xõ�f%��9�b�E�7�AO�"�\߫��[��W�C�}B�}�Fj)*'4��k���ef��a����@�|��9����L�dj�p�=y� �Q����.���v�i�Z����~�g��2ψ_�~L�?�TzM�f�PEz��!Q�b�8�Hcǐx�;|�XI:�P9��D��O����*�t������D�;j�q�|�?�*g�F�ECH�������pN�8�y�Uh!�*�tJn�<� ��%{Ԙ���P��>n"��@�� ��شA�r@��Ϛ2�=
��qd���u�BR�M��Hw��.��e�"�u/�V�/�2Y������৿�F�=��L�|��\Zģ��[�Z��K0�A�7�`��ׁ��>Y��������DI����*b��@w#S+������@%c\7��m&7���oء�h�z8��Hj6��dP4�^ޣ�7�E˃,.b���^I�?g��s�"JR�2q�h�xUY�w��c�w���&�
�O�ߩ�7؄!��!p�i���&�#K��ԧ�*�Z5�ոXiG��;@� �d��<�V�o���o�R�M�b:�#����q�F�1Nԝ4l<[�N�Q^�$��F�g>t���/E�>�j�a�XD�a�F�AX�jN���rH��&�<�%�>���;�R�5&Pކ&^�]�)�)����5�)���l��	�L���P u�$n�g����F�q����e�F8r�����P^��FŻ�/���h],�Ԅ��75
�ZWwV(p䨱��?��1(Gkh�yL�@��Wj���G2�6uG�ǉ�"ס��2�Bۍ��+س"M`5�Ju��;� �1ϼ����,�Z5j��lڪ��9^�s��3%%��a�c�і�\�a��R9�^�ٺ3tw�CH?�,���]=�� �B:��"@��-סeん�-c�/��޲�����K߀nj��y��H��T� ��.p|�������|�c����%��
ۙ��X$�6.@��[�e{0��#
#�[�ΐ�H�r8^޸�����B�,�g�o�\��.	�j��@�ko��XGy�f.��P��F��Fn�G�7���oߨ�]y�R?�M��m�	�%�(b�i���I h��~:��"��%}p��
w�z���gY�rG,#F � �X����i��$"/>C�ޟ���A�����Bc۾<}I_"�gz�7qh������]#7�q�'�rl?��ݘ-,ob))�.�d�8�]�.�yK�c�4��LA�L��}��%��=2�s'ÅPH��سy�4RΟ캟�!�9�_|ٍ������M�ż�t��-J�~fhI�x&A�/��&'ބJb(��Xn�Y���ޥ-�6)���2�9 n��|��~b�Gb��/����'��+/L�ނ���qtFS]���g�%v|��K������g�!T~홲��L� ��'b��f����F0X8��ZԞ�/��Q)��)H���Di\�LM�gr�[���p�5�J�w{��1~2�υ/B�,� mI
"VË��PƵ{��d�iF[�BK�����_�*�5[�+��g���$�mD�ʢ�K"[� d�zbQ���kkI�����)}��2Fr]��ބ�Jm�,(S�0��F�l�a�	��Pb���Yu���}aCª�(���n��oàa����)���mȥ��d��c���7Z�S)MQ:}��J������m��v�.�,!��9��ݷ�-��Z��Q��UP�J��԰�IU�5��u+Z�_����Y���H���oD���`�I�/����܏�i#R({�B�\�M�JJ���,8l��c⺼2�(2�2�����(+�S4/�A}\����8�*�߰8U,�yU�z��?�2q@ �[�̪x�g�v]lv�����j���_vZߴe�}*]��+�O�%��zd>��ᢀU}��%��[�g�4~rID<���ӱ�S��>k�ۉOvk��wH��"���pa;��5׍Vc�QT��
��L�����"X��)���5��RM��Y�~.<g�5����z�3�J����*$�U�V�o����J�?҇s�8�a�$�1?�NO/?:�f1�H4�k��ܗph��6�GQ(x�H	���&���*f+�g�ki��IR�{v��I�_��c�t�h��|�dn6��~[��6�މy��ts7�3Bk[���A$ǪS��&6���B_d��<��^=��	_Hߍ�E���_����~�o��ݭ�l�MZ5�c;0��t>h����Ov4�������m�*>�Q4ʣd��G�pyS7�Wώ�#~����\ʮ�� {3�
w�	��)v��	$�Hho��W��ݡ]�|��{��e�$�`�����tk�B��s^���Q�!,���ۂUw��h���S�#'��AdQ;GU ͔�w^���t�Hm�L�o`k-k��Z*�740���}�k����?hF{�	�*~}	՛s��y^9��⃦���#��a��tʲ, |��X[�Y�i�}��v����x�A�Q��]�]�� ��0`N
V���w��ds�B���L@��~�QY�	b������q~1���z�5w�z3�U�W��>�� }g{���prP>��=Sg/fR�k0#pQ����뺒uh�u�E���;��rvd��>��jm2�\6N'�%{��mg>\��=Z�ݪ� n[�1Q�R�Dq����2rn��4z㋠M{Z�ܚ/	3��}:����|7�:�}A�aq�����efXU$���/���<� �����c�_��sSŭ��4IF�������x�Z�zx||zˤ�#���/�$�;f׫ �D�ͳ	�+�A��_f@4�0�I�'��[�}��r�dV*�w�Ƈ��Ѿtز��Ň�ɟ�X���������ʱ2��䕞�MY�Z��ܕY�9��u�_��R��˩y �'C�࿡�Mr�My���:����Ã�рKV �R�6�ؐ�܂�T
*bV�,:A���u����e-���lG¥D��NZ���� vfbLnS7TQ;�Ds�k�\d���47?|���ԮxB�ۜ�_,&C����v�
7�0m�=[��������ͨ:[;�}P���>�"(<
9Q���5�gP�Bш�6�$>�S�����ډ-��P������Ӣ��A6�|@}�)�����&�E���Ԍ�����+�:-&���:�L(��@/S�%\�s���x//"�X
BZZ¢�����A����>���
������;X:�~��K�bS�G�w�)_Z<�UoFs{��Bn�����?���Y�9��O����«N�y���
<u�bVQ���\I�PU��i���Κ�8�G8��E"!�D�ɉ�W�~�Wr�.�����?�)���1]-.�L�� W(��T�����9��`B��ށDʝ��ב��8�����8��f��d�A�j��c_cL���FZ(����3&J��;I���j0�Q3D�R��-�u�&Y�Aꃨ�>rH���E �@�EN���J���RbG�M��+�T������C �5����:A��*�^u+]ۿ�������Z�1Vdu���Ck��<�������L%�5��j�t0�%�|�`[����������?�gQ��Z��b��G�(�{U~�+	���o���9t��U�N��x���_�ue�.k5�>V��z�+}�5�
�!����&o��^�Z�J�2�{B�>�������*�F�0s�����-ziT^�����<N٣=��B�< 5N�H�wv!!P��~2W	�|Vq�zo��	�r��3��	��sI�Kc�I�C�Y״ș�|m�cDj�6{P<5�&�Smi.g�ާՀ7�/O���eXG75f��c���6�^ȡ,i,��h(2H��z��"n��_/~�Vs���L�,�ꃝ-�q+J߄�y�~/�Q+��Er�F����y}J	\��	�PX�`��#p/7I<10��0<��a�'��k���LA�~�+��_O����e���$��O%�&����,� y��&��=*�Ln��x�!&��I'�.����|��07jf�뙍�hy�Y�GF~Ua kGʘ�I�E�U�ou�6��.����:�.�c���v\��(w*\��"�`J)��5�����@���{�|�O��d �(븍�������f,�f;��D�b�>xD"�P�{<:v����eI�G�p���`FQ�?V�$|k���$�����RK�j����	��������%S�}��߇a����"����6g���Z��|�c��BK�V�
J�/b!�<ԗKӗry{�hH��~�4�5�����^��LX��[yv������p0p���
:-��ؕW���8����a��N�1�e8�V2sQ���҉�����'���x�g"M60dt��>�v��ᆟ��?p��{�Yw%��o��c@�$��������m:��D�^sW(C���1�?Ԁe��Q&p�FށۙID�IG��`��WG�4�P�G�]���#����>����*M	ϯ�L�K
?+��#��&�E"6Z��{�:+�r,�9��ֽ���C# ��^%I�s��ܭ���2���x�3��6�h{���]����bҷ�(ʀJe��+n��Nw<Dx"ا8&	����8�B��O���$�H��Sf����<��_�&���v�wd_.W��4m;���TE���W�-��)���UA%1���,��jBO^χA���������|d&�j��8�`�|���� ��-���h�����pA�~_f5�G�Kv�s��)�H"�Qٕ�L)���Y9��p)���n�s��=y�ӼR`^-�V��Y
��4Ņ���
���-FdE$mo%��Z%�j��\�`4]�qd}[��H��4Va,��Ƣ���
ҽ$TdB&�^��p�n}<;�T<�d�"jo�Ǯ�^RQ3ic޳��%�r�b=ɱAm�r-��DL�B��W%Z�驺�dud���վ7�qfwAk
�0VO1��/N,�_�d�2��� Huc��3{ÿh� ���b�����wL�]FU�8��%�����<X�^"_��F
�X0;�Y;��0�K���Խ�ԛ�ܪ�"��Ͻ�rgu�-�?����!�4��&�W���z�Q�m]�Ne���Y�c�����7�@A�v�����_{Ҕ9���P��hd�hV^}P�Pb��(�w7痿��d���[��CҨ�� �̡��S�~����t+���5f��UL013禵��������v3�
��M#�+li��5��YW��� L
�2S�M�P'��(�$	@�]�9{���poF�a5	��#���?�exj��Fd��^���yF?[�	����' ߍ���#lv�vw2�, 0^�v&��2��?�����:l\�Z�G�.�-�^C��M|���kQ!#��i��װN����������H���D�}6]��`q�pG����9AH�Ww���2N3C�)��W5-��ʐz5��ߚ�pl�Y�L�h�Eț
������(�/�=%o�9kv��޷� �n�,+$���Y�����������3�<�C$�7!�U����� 
�|G�z5���[�Ҵ��87P�	��]4'�6��cBq��t�g�W|��s��=Kk.A=�=m���ȳ����G����_Rq?S	��_V�u�����Eŧ�չW#o'ӏ	�pj�b�V�@�/��#�P����8K�)�Z���N�Gw�2Ueڤ�5���l�i����At�������r�$�Ҩ���;|���҅oSG3n۱�'SX�b�q��)���Ic��>{�Z �k�#*ͨ3l�Ǐ(�K�ch���E�ص1���:ޢL��(���5p m�����v��p�K�
|�+��������E�̎	�n�N�@��]Cl�֢�eE��[R
�~�}`~���hp�y:X�u{�J��{���Y�.Dx*	�j�?�o�~p��?�*�@�<%DAw��)��3q ���HOvI�jr>m�s߾�KF5b��ĆJ���G� ¡{C(L\��b����x�7�������lĘ�ջ�ՊgL2_� �������N���-�&\H�`�Q��4RZ=a�d���^��[���&%Ե���)�������@��|��O�$趒�'5*<���i���>=k���Dk'|VI"(F�F|��\O���G2�5���į�K����C��&R���x�(΢���)�[�I��t�uBϐu-bW
�v��jt;��x��ݚ#�ٽ�YssQ��Lc�š슉��d�J􁖷A��n�H*��0�UC?6.5��Y��2OK�?��v�E5��6�c0煬޺�9�$r��lg|�ۮ��$M�����D�tI1��v�%�/��J�-�5�4�c{�N��8�#��.C�Gb�O+M0P���ޓPac������d���v��p�h6���%a�M7�j6���c���J��2��|�[����i�"�x��ƌ
i��5��_��Z��ŧM�U�C/fh���|as��\�{���k<DqdUk<��>�n�'�$�H�Kx!�A�!���L�3��h�����9XV�l��ſ�"s6�҄n����sD���>�ܮp�����B|��Q>+oI{�� Kh���`��K�`
���_��[�v�_Fŭ�h�־�ds[�X�8�<�a�!?����o:���W�m��E�r�!��vJY�~�Hq[�ַ �)W��{?F@#�<��'��J���*�ā�};D��r��"��>�<�Wr�?X��̓ldۓ�=�Z�
��`��'�cN"�̄V���tO���Q$5	��_J��I`��_J-�?���T9�1���vf𦺠�.��k�ـ�_d��@^O(Ͽ�oLx��o��� P�YoJ4��BZνdXiʧ�,�:{-49a\����X�E9~�\����m�td�$W���MO�I2.q���M�p�����6��#�uY���m3��xn���vC�)�MB��n�Z����$b(X�{zP�h���7XͰA�JX��P��Jq�_��:C���;�G{�^"��[����O��Ӛ��$�S��0o�5�#�|�Ѐ��IX��oS�^mp[������C���/F|R��S�AΈ�2�e�U�'>��q|�����U^���^�r����O���߯L�nP������%jݔ�i���(��*�2B��c��B������/�S���	Q���+�e�а&���]ݻ���#��$>��mb����V��Y`��=�}�߈Z�&uMR��I<)����C��2h��k����\g��J��4���?ֹ+jv4��h�Ib�v=!Ĺ[�m	{��a�YL)˚�"�936ǙI]&̪Y R��n9�������ԋ����|��kD�d�ܯQ���)ܛ���Uȑ	lJb�Le�u!��<�2�_�N��t�����b/��wlC��ϿrE�s�rY���6�e���ID��mz����=҇��댩+Ke����;B�aΙ^��r��`BL�M�톮�V~ ��, �q�/�Ck���^��d(��N��¯<=y����He�)�yS�W�A�<���D��	_�xi����@�Z:��,7�$�.�	�r\��k���v�i���h)���9N�-8���2��i��.;]q*��X�(Mm*0e�Mŏ�/Z��EO�gs�	;ฤt#�Ӣ ����[�}}~D���Y3�6˸<-Psb�k�����c�`��?C3ᝓ;/�,�	�s!�g���oE\�1�wmv���o��7P��	q�
CDxi.�&���"چ˲S G�p]�9��Lq#�~aWܸDBe�n��������C �z̍"�3��8U�DkE��x��u
xijQ�e��?˔H��mM2�:�6�w���7��⪹��ҷzl�1#��7$&�7��*'�����CP���V�?����E>�V\02�Ǿ��Hu畂+]�ޑ>RS�IJ-l�Z����#��}*�KcW�kazb�h5�Χ��|c< ���Q�-w[<m�$e�����~L����U�>e�]�˕�Y*+�s��N�9P=��U��Q����g�2��I( �i�ɛm����p�hqz�*��e�^-\���������❩��(=/��L�ָ7�iin�_&'��8���]��3a;S�
�ݗ�{>>���e�nAj� ��==g��1�eh��.�5��v����UX��6�?j�aZ��QAnVB`�+s�̜��`K]�<����"����[�찵���^����V_�%�58%I�%i�?ۛ��:�D���m��)�2���� #,ue���Ɠ�t�S�R�Ȫ��@6ƅUs��ZV	˴���b����R�8D}&�X��|u��M~m��F&=�+9�Lk� �)E�ϲ����nՎ�9q��25��
Cɱ}Z�M"����xWV�ؽ�7�)y�V
�� �Ȼ5���o��.#�.�8�֘k��d�t�o���v��-�b���iu������+x��Y{�L��34��"���8�T�H|��g8/Cq/�U�����K>�C٠v��_�ݓ��N��_Q�~xc^K������Jk������I���l���>U�ŮpuM��h��:̚t ��|\I@z�ub������@$��w�=^~Ѷo��^�7�c�-K��W?M��������F�_�#j-�G8��C�&P$��f���a.w_�|�c��5�aT+\$�K�F^+,5l&<"x�9�����v���P8){�[��#࢈�I
N�V�o��H&[/����ߏd��� t��צ9(��-�����/+�����M��ֈWi�4#�Qw�ʣ�4�q��u_��W���ֈ9�h�e:��w�����'L��k�E��*+����RM+nQ�
U�ς])�<�ض��w,�M_�&��$ۘT{�w����B%ی��;�2�7��&ixA��~7¬o=��U~`���G�+[�Ǫ�)��4h�Ph_*�[�қ�x�n����Qƞ�@n�`�:D7G{�x������E��+�J�R[������P=f^ݤ��	���Fd�!ɟT��o;�>.B�ڧ��{<�9|v��T+���G���lǺ��=���#��k̦��\���C!��A�,�T: G���|�e�y�{V)y�(�J��!��@eb�u�Ԟϗ����1uQ]
�1�˶{��bGЏ�)D����?[�*��T��$��� ������R�淍���P7�z�w�S�-c	�U��k��=}��л���*�\G-Q,K������ ���7���l� �%�K�V �Vf�Ѳ-�'P�g�3�d��;Ҫx�����,Iy$���eT��0r�&����I�sӣ�A;��wqy"�=�]/���Eƅ��_�i���_8�����÷����% ��>�)n<�3���7�}%I�A�+�^hQ/B[�G3�:O-Yi�"�f�?{�p�q$�^@J�gn)$jk;?���@�.^#J�U����f�_\6����H@�2�ͽĮ�k�DͰ�$�P�f}����d�c�6�(���r|BtB#�	%{�B��������-~�QS�`�J]d�/�â�*��A�O���I �edm�l�#6 ?�9|0�O4�ٕ*��\O�(���h>@��z�E�Ѩy;x4�l��ҝ�b��[�,�\��v�9�Yd�������Z|��i��l1zo��c�1X��pŤl4X!���T1F�v5�%����%7��U9��^�J�	�D9��F#P	��>8R�FS6���S�l�B+�t6.U3����N�B�K\&���C���Q0XX.�R��Q�J�-�z�E���9��|�����o�m��tq7�6#^�	�����4U����x�^�\��ɮY�܉�:�E���M(G��0�1�J�=���$	���sݶ1ю�ܤ9��]k�c_ �]���SJ����`/۬f)v�"l����j{���P�n�������!�]��w���\%di�7��� m$붡95�.ǵN����ѰI��K��<QB���� �m��r��.��A#��Md�k+D�3J����T��H0za�:6��L}URlܞ�	ML�����==7�o!���' � i4��^��4DA��}(���U���i��H��rm�:t������ʖ��*4
��ȷ# ���L�X�D/8<r��#�b��De�1��
iV�Q;/��lY��%ʎ2vX����+oy��r;�EǊֽ!)��tw�%E��J�.��^:��!�[��~G��O����R�_�)���-"����,٘B�����xɧ
�*]��8�٣�|
�#��C�]��32}SWMkyzJ��Yz�P���NM�>�.�p���Y%o�A�oɤ�(�p���[g0�x4⺩N���
'z������s3T:�Oi��,��)��YsK��*��Mk(���z�u͚��=���Y'�5��]Ӳ%j��<�����QK�G�+���v��tB�͐oa>K�I��O��P�5��Y�Nk���e�܄����I��:T�S�<���@u��G&1���B}~)+�B����>�\�*}�5m�$��Cx_f>.b��+6�Z���lS���z=l�ZX���3C���U���,�"�Z���mz�;ƃѾL}9#�x1/�؜��(Ѐ�zȑ���$`0-�ǂ��O��`�����A�T��+��)���0so
�#0�lX�W�P5+9�N��ˁ��\� ����a�}0�7�j�������f��o�Ss�/\�Im5%K��z���K។���j5�vB�|e�m���Y�B�նd��,*�ߺ �����S\yŸd�ŉ��L����T�9~A�خlҹ.ݖ-3Q��)�~dr��z���Ү�����_��Ҟ�O$�$n�:Oɚ�_է!jjc����~���o� �\bW�}���0x.�u��,Ѡ��5��%ʛ��u��ù��:_ǳe\��7ր�Y`����8y$ª�`�L��cl󝀳���"(] w���$����H��i7o�fɠlX����G�U3c%gO��V
M�-{�׸PV���<�5ш�~86���\R�X�w]�%7�0<���&@8���"��fڂ����m��x|��tU�f~�x�$ޗ�Œf��{���Α�u��d�;�9�Bxh�����J��G�V��c ����v���s�������N<y�����b�n�y8W�ZfV;��E���$�Z2�j��z��?뻶�E�
oO�h��re�[�$���y!+� �j���.���S�Uj7�)~�v��
�ⅿB�A���]�CH��&�ЬDJ�Ŧ;Lp�Z�`���U�v�ט�=�!�I;��s�yO�>�j &�9�&$ʸb���h����{���P�@-�V��q͡���cG.1!s�`�Ƶ����Я�p���}2�k��B;���	%F/��'ߣ�qf�y��y����4���g1:g�V��:�]��߅��ٽ�#������S�r�}��2 !�َj�_�6 �,�w2E��Fs� F�}JC�O�k�{sr��g��%��H;h�	���)��XtV��S�����#�-�^3���{^��w
��h�ݢu���9;/�>u�#a՘���9�*�c�P��������S
�B�V3߀%R���K��_w�_ ~��\��`���
Z���7�B�ɤˠqx����SD`������J�c�{֔��]ձ:("�kZRU��:AW��J��_%�M�F��]?T�(5v>���)z��J��ڤ����b�u�i��Q,i�
�n1�;CӃ�R ��hξ�rkR��A�����j�fqY_ڊ.�e�`�S�x��W�؝�M(m����J���ݣ��%�[�rA����%bc��k�?�4�V��6��'~�o��-:1I߸@8BMG�e��F��Y+���㎵�cxWO\e��'/ ��o�C2x��Nڌc=��j���¡�0�b-�Q��:O��N׽R+�v�j*E� �?�G��/YZ;��&o�i� 3��EQ��������7x}ML���� �>W�A�#u"��)�)���d���F��mz���˝�=�ބi�4�|_}̓�1����&ݘ͌y������t?)$�̕�����2[x���S��hb8] ��<a�����e*���P�H��˹�g�E���ٺJ��D�v����S�_(���e1�z����=�^��pHQ�e͞(KN�s��zJS�M��Y��L�L� hT��m,/V�n�E�)�?L�뉸�"�z�����*)X=]'qY�~(f�=�4(�.� )�j��¹��1�nt��:��aK�,Е����Z|D��m|��G��1�V[�&�/n���|����tQ��yU�u��$�+����
T4ܻ��I�;����{��� Gj�嶰��]8�k_P�����94�Ev']�P��Jch��� ��,�V�tB0�;��u�B,O�A��
����FOL>k�z{-���'�:�o�4�H>YE�]��m����j����xQ4�Nq�ۤ�DP@C��N\���^h���m,[��#�p�c� !2�p��jYBf�7��T���*��Cǵv��7�_�@�����KE�KM�l�d\-��6�l���R��[o�H�IҌz���ߖ���nxc�Hj�3�H�����؃JY��͡��5r]GN:Rl�qG-�h��}m�6#�3�S=��=̻ۣ���{�������݉��LKS���b��71)y� �=c�JX(.Gԯjl�ׂ����b����Gh ��Q;>�q%�K���`x���Q�gN��"��r�'�$��~@1%�eIjɎ2�ToFU�~����T:��X��i B2U� �vO���i@�q�(�����4����w~)׭��a����A�{����o�\���C�h�a��x9ڞ��8@�F��v�E�I�gN�Y�u�X���&��H�E�}�2��+�-UGg�,��� ����&x�a��XEHs����M���X������g�ܽ�Lؠ�?�A�@g䵨�ǀ�2b��`��fd���H<:��̬�N���V{&�y&�N��+q9Ƽۄ�w
j]	����Y��r�#���;�}�T��l��hn�6���FF��6'��,�!O��%��g�|"|�Z��q�ܺ�u�ON[Cc���!>��<B�K&}��9Ņ��b�?�3�N�:��u��/nFz�h�|x��Y�`�ts�+��MU�C�x���:y_�����aLe�XX,W㨨q�A��N���3�����mj����G���P���rU��al�U��(�µ��nL]e�|�[�$��E )���R]��
�c�:��C�X�`7<�c�>q��	:��] �p��#S���:�М`���V��y87��������dBӽ�*�z�k�>�ۀ̷��|�=:������cB��7�%�a�Ӿ��g�e�����ז�Y��2�v`"ҽO�t�g��g�N�
��1��x"M������k(��	n=�$L�9E��)+��5�<��E �)�$	>8a����^�L���	����)*Ul�1��].��z �D��I�P\)�E;Uך�T�p�����Po�}���N��b�m9�٫�J+�Gn���!2�«�F��󀠱�C��o�P	=��i����;ÿ�&X�8���`n�ߌ�TŹr䷇/��]�%�䒞�1|Љ��^"����[�1������7:�����1c��:�z��.�cŰ���]�O��q�:�6p�{&=B�Ƣ(�����C�U+�P�'�0�V����o~����f�@E��^8"e`#<��J�^A���m���z`	�VUgg'���{�1����y�K.Y��A�������C|�x���-F�%� �o��?��Ls���Q)�9}`����P:��+@��VM\�Kel�lh̰�PX�CK��+�5��,֟��N��;Y�ɸ�x/�S{�3
�����ؾ�t��T�n-�&��:����w�F��<�������Ԉ�ZH�+tz��@� *a��j��!��;Ўj$I�+0�%����C�Q��8W�s��$���&���aX<����}y���VW����U^�B���9EFK���6�����cTc�)��׵ϝ��[1��ߴT���@�7��<䝂7��c["����O���:�G��#P�|�,$Q잞�(�:tF����m��bP�6Z\��q�R�1C�klp��\��[k�B{m3z���ce9'_�͐�&Nil|}a����'I�% �b��o�����n�
�ݰb��i���w��j�]���`�:,�X�w��8/n���or&?|�g�Ǿ&;8�F��t�s>*������6_W�0e�"�ܜ[�rl��	��������A�ǔ;K������r���U�-�-;��?]�����;���mox��8R�����r�s�DH��:�}k���H���ng��Wa�A�j����8JC�bT�6��.�JXF��-�0���Y��.w��B�qȸ�����D��^ӫGl�2�f����Qi�u
za{	o0�v	ˡ׬&���ȫ�<}��Wl�/�L�b4`w�W�I� ��)�VZ35���{���^�ݪ�ۼln%�C��CZ�|Һ�9;lOvw�������V�gg*I�֑��G.[K�� *b}wX�����+� �;f��$�yy]�,{QU�9�=�5�Ǻiŕ7���Uem����_y��ܝ�!� P��/o@����ʽ�����)�vZ#}\Nzt���7�O�ǀ<���[q��2�	D�ԧ49p�mTV�w9R���9�(��_�B�F��6���o��GN�|���^綢 a�g���S�[��$���p+&y�3ny�^mgÆ�S�J�.��x�Ph��o�^��Ɔ�*���N9 ~Ϯ�ڌ*���������'�)�`��شo)Z���/���������c��B&��q���֏g�ԕ�Թ��ݵ�ɚ�^m��u火�x�=U���W�BI?�!>�@s���:ʓ���9�3��	�?��y���ȹB�f �(y�g��q��Wg�@�FXI�y�8�q����+�/�@<4k5��`g��f(��k������ !�ญ��-v���X��X�ɜ��{��	v�td!v�p̢�#�&�ӟ��+%U=[Ę\P¦[$<��4����AP]ތ�G��>8OR���ߥ�դ��O�2N�K\��q��g�9o�(�8ҠO=��C�2-s�Kv�F��zxWw3F��%�řk�].��t��]�!-�m-������5�����:D#ݐ���B"d��o��&O�Q���
-��M�k�/�D/�"7��}!��\��k�" �?�m�B�3��y�%0.�p'>�P��f��W�ۂ�ɨ���pGގ�c�C��g�������0��T��7ۡ�-�D]JaT)m��'��]���h��m�J�K�FD�J��* ��-M����N���~�ѫ�:ф������?.Mſ�`�sECS B��5"��Y9�۴)�$ $�V-����d lN�Jtĳ.�ʇ_ŽNIx���æ�|E����4C���y�!rcb�k2K���7�u�<�݉��m9Ci��8�9O2w#Y#w?�Ł�򵧍�g�+J����w"Hɓ���(�x(9�1�E��Ɇ��\�#�F9�&��� V:�p�W��~rʃ?^A��,U��TkEÁ������,�V����a体��(�)'��q����j������7�Bsس��ï6�b~��am���J���o�LS{�ag�����Y~�=q��;5U�vzox�����W�M�����jn�c�+���l_.֪"�	f���3Qa[}&�sϽJbߑ1�z,Λ=x�� ���>h�ҧr-��w��� KT��ʎ� ���Kl#���W()q0	��σ0��W񫬛�%�~"T�i1as�}&�3�a�@���B���jQi!
w���A����_��6c��ҏ�� �>�T������R#�Zħ�w��jWZb�1�	��oA��k]�O�d�anK�϶=�Ďס�b^Ȃ`��[�� ;�+�8�]a�,��5L~Aa��lS��J:p`<��|`f�Q=[t���hvW3�X�P������z�%0@0�R�p8��}p�����~��r���1�5��E2��5(�����d��.]&�c~y�T�:Ș�����J}Uj��#�>==.gj3&J�I�:~���Uq��.y{n�����ܖ�gů�
�Ĳ(f� �lB���뜇r]%@[MO?#�Qxx�	�`��	rZ	�{�M
E��HC�3�N�#7�"���p�/��c""�Ok�r�<�W�1�_p���~���^o��uݜ�M0���qჄ�[����OAnk�?���T\{�mV�V�wyb�<��$�.&�Ӳ/(5E4YJ�!�l�u(��d~C����9ߩ�V1گ�R��}t���w���:��/�t�
��v�Mʡ�y�8v �Xt��N�~���h4��('*C�:o$f��d7s~�]�Lx�tAZ,��Q%��&����B7�?wb=�S���qx��ei2�I]�4��PB2a�A�6���\��6����s^o���g�À�4P���oH�$B���S����mn�7b�;Z$aqb���Z��1 ΅���U/��^�
p���� ��.C�l�&E��l0��� �N����dw�oe�9�i#������$p�)�BV�PHg���}� �ر뛛�n�B�����b�^]}����֚̃ĔT���u���ZO��ۮ=<Q9|���-	���X:P6/���nb�����\��/$$9�+�����.P�t�B�R���[t�yh� 3*�r`�)Z)��O0�ˌ��Hn������V>Pg����-D=�*���-��Z��^u?�^=�P�����͍� R��ѽ��S%6g�ǁL~m�+N�a��$\��'��ؐu�H��'&�F;�=O��oRP���6lb<�d9Y��l����B���+����)�q�P�l��yGF$L�_7s{p�	 f]��F�vb�4�����)�	=��r7%O�8X�ّ׆͞9|���GS�f�Y	e����Az�i�O�4��rH�����8F�����uG /�ؼM\v~�Ԗ&�$��p�4l�-�=�}��9O-�6�>��%K_���&������|+tj��y�Z�)#6�WV0)�uG�K�NE� ׊v��~l[��m)�n���N1~�R�Ҷ�<4@�V�#g��V��o����F@q�l2,蜶��3N��[��|��Ǻ�3>�W:��4:-|XA����ٽH�S�ȫ���^�˞w*�Ä�IY:/��9�