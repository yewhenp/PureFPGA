��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�/�E|$� R����q�m)9)�L�@@���>�@��#�φ�i���wk�S���+�ADW��<iw��y��+lT��d�Y�����"߼�a�V�O�)�g E���5�e���U�� uxB
�;����]�#l�'x��#��A��0x��_u
ӫ�����(����J�12�����
H���`���"���n���f��< ���� qz̍��Y]<��wɴ�Q�&�|1Y'f%;�8�޼�6<P���x�E�礑��`�i��p��o���4�pRt���T�V21��n�|��?ݺ�o�3	����!�F������S��G�����3S�=y��_I6�T����*əA����	"0����冧'��{9� "��둊W��㸧fu�{3k��^��N���0�3�w-]mM����C�h�4p�C�&�����^�ӨUŏG��6��̀4�� o�!?e�by�y�����c�j8��1���ĩ=�jnHEx�~oYm#d�w�wh�B�j�z.���O�����������bQ �*Od+6�q�E��P�p��%�v ���4�D|��Q�+���>h�|�'R��à$}��q�,m'i�H��`��|�+�*���Vv��Ir�&�`p�;��qg���n�a�J����t�U�am�5	�Ϻa%����۾��{�4P��\�9`��J��&񵂸�qzfV�J���^X���?�?�pp�APK)�:�6����gB�E�F�J�����R7��C��y��
W���ƶ#���ybUd�I�F|=�L��������ld��^/4�>�IT�J]:�/&z�u���^<gֽF��Vok�<ɰ(��6޺R����\��|�G�`����NƱ^&-5.��PZ�Əbo׽MQ)t=������L�;�f�*7 �Q�|��/�n�?�h�o��l�����;���#��"'��;)	�p)@�3���&�dm�#'^��l�=�|� 0��u��uR-���+�]6K���^��Q���̾����	��fR�Ú���NN�*L�퓣x"�%l7%Ü��Ydx�VNK��aSӜ7����߲'/��������O~]uE9���i�uIiʱ����w�*kn�y���2�d��n�.?��d��y��ݫf�L{�s�����֑?�ʄ������A���<��]�/�@�A����?�Y�]������	y�8!�.���]7�@��E�B?F�I*FE�]9�8�����V!x�,�V�T+:=����3��#�p�&�0��f�Ⱥ��?z؈�4>7�ʥ�����(�J�w�l���SM����n���VḦ@�KA�%k�fp�sĮ��z��5���O�R�N�,���HS�S)�8��'�}�"T�9�E��Z�Sm�!Ŋp���7h^6�@������S=۷0\@�xs���ǂ�`���c	R�/��a����'�>�P؇Q	�bD�M�k�t��s�|�(6�y�ȉ�'U��_�x�L��gFF+��}`���T�u�����K5�Tr?���g�G�� qd�Q�4V�u.�ѡbѿ��ʓ���t"o��*lF��R��y�A�`nE9�<��_G�FQM�S�К��~'t\��|�z�$���(�i��W��f���~��q#�����#KW&��v?3�����[o�!����dn���@��?nWf�򹻬��y.�OL���A|���v�Z��X�s��؝c~NJFR8輀S��G*G�)eL"eïs3 h�X
E^6\r_�!m���F�nɣqA����,��BT����;6u�i#j���R5ɽCS��'�vS�����V��S:��P�l��H�z�<��>�I.���O��Vj�������.])P��X~���D�$�08dv����,���9�6�i��;�-��+�M� �O�Am�3֦��r�nOA�?f5\�B<�0C��z�&g�8哰xDuJ�����do�s�6�h�~|�%���P҇ouZ�ؒ�H�>ܤ�c�nqn��E��e�%9��h�i{�M*hO1.�%�,s臟�����;ע���sS@��*���y+l�g��i�~`g��I���TU�a�$�
 �D*,����8g���_�/����8��kX�?oڳאc���Yb[��<��Fݟ�J"��M�r0��zA��CYVs0ꘁ
�o�ڟ�t]��[�\�rj@���2���n%ז�؇LB�͌
���kEܼ{0O/J�**�z&|U�f0�_��R:��T����gs��!�.�;�fg`)~�ƃ�3SJ� ���x���n$�Oq�EB��Ն^��8�$��\b�[q�(;������t{�1&�o#�2����@��;� 5��X���'DN�YZ���~]�:f5 l>�nz=)�j��jl���6�N �j��9?�����	KO��X�р�Fd��m���r>��V���g°�K�m��&�&�U��.���DK�h��t��<�������h�Ů�0	9��B�Nj�ٞ��������߶��r��\��f�S$Ƌ/SӼ�o��|NjE�xT�O���&����[�Tu��܁dK�H�T⽪ˮk�QrD�Wp�iH�=�G��H����N���A�z���'��'^{���r�t��E����IcH�O]�d���x-e:���F_�x�[	C .�
Y�}��iu���(ψ�)��Mj.^�jk����H�~J�x�ș�!2-��pf�8.�8R���s_s�	�xZ�qMM���ױ%@�n�42�)n��ЃI�|g���X���O�בt�sЍ5ӷOB\��ԣ�]��#��0{>���e����BN�����+{R��ğ�1��O�Bׂ�t�}@m������/�P���-�d�`f�'���26P��~���+�h^�������������ġ#xyw�.�w]��u֋�ѣ��y����YYjM}�D4w��kؖ�9��ع|�hPu��,�&p1n+���'��̼Q?��t���Q	�%��KL�b�V���Fvbf��ps�/����z����ҽP�������,L�&��ɓ|�;�guى�;��~r!ZX�H��/��+|G�������_)�g�����v��й��6��ڛ��_؊���@��'*8�S:��G�A~^`�A�&�7Z@E^ײ�X^>�&.��M�K�o���Z��>H~���q��!,���
B"��X������R�3G+#X,��>6���$�So`;�0K�,�|�nǋ
��1df�',�]	�� ��MsT�M` �^�{^�+,<���q2�"�D� �ww�| �H3�u���
a֎��6Ĵ�}cp�T�U�ِ��X6�8�����+�ο��j.��H4=z�N��~
W.��j��v-5T�6�؀k�}�~�3*�WS�a�P2�����_AyX��H�doݽ�ܜ�M��Nr�.��?��
�[쯵2����m٠�#�yV���GIi��"�)�8��YF8�.���A�U*u�I��n���NzzBG��}���q����7��"u�>���n&ZZl-�/����WG��AY����p�Ka��4�nܣh�h�D�f�
��V�7MEz�\�&4Ç_�í�+`SA=��.׽��{2�DD��J��SPǭ�_�ohR���}BL����}���A��ڇ���kG9����a��{j6-)�/��#��Of�x��u�JZ�#d�az���=-~f�k�"d���)����p��f�/w�� <B�����R ���ٹߦ`+P��*?������m!�fEy�x	e�G%�ӻdE�G���=4X?_����:�?Ƹ��e"�f�DZd�Y��Z�o��V��H�<��na�r�ykq�T�'��IidF�e2��NU���=�*�4�Mz�'���3�М���ñ�3�a���_{-,�p���yP���#í�DB��D|�]Qv�.� �Y��9^���'�*��Ҍ)9�4kh4�g:����\���>�u��Ѫq������$(�;�D�Jb}����Sc
�|��y�U�3'���6փbںyS�s_���necUs>O�3r�0��d�OPJ<B���T��k��	}�u�C�f���
NX��\�cw݊x�}i�\����z �'���7fZ��J`��,�r}2�E��3?`���󻈯�^{����/���d�=k��J�~u8�î�o��އN�	]��H'�~� mVD��5C��o7��v�U������ٞy����<Rg���NGݥU�����b`(��'�����Qh�V�߃	y�Bs[�8��C<\��J��NЪK&�g6�)�|�`����W[bp�M�k�t��<�`�QW!@�̽>AK���8yF:�'_�i菛�)���:r�����`K'�bSɯB�Gf��ڷ F*�е�o�%/A.�0��8ۨ�4��zL:�5��Cʴ@��+�ʕmJ��VW
YBEZ�>c����I�9���9R�Q��.���fw:y"Q��_H�w/N�k�����ڦ�&d��wfi�
�;�L�����	x�)�8���"��rX��{�B9�|Ɂ.�y����wȮ�_��<s�'��+���6)�������l��qS�<��e�ټ�{"TĢ��c���HH��� *���Ӗ{�I�':���"���C��Q�8�C~|l�x�FOi��aß��R�v\��ۤ'n��慵��"��v)튑yK�,:�/�R������=��ퟶ��Kԍ�l��Tͪa�r%��1��4.u�T�E"��~�u�V[��gC��.3�X���)�Nw���96h9ޕvb�˵�.y�AZ1����il���.��3d M�Z�T�0d5�4��
O�`��ʼ'!���;�>	:�OEe6N�C����aQ"_Ĵ����rc��@�o�����d'H�����g/��P�zxRLz0++���C�~z�fk`{�O�K7�"&uk�9�b�:"��d<,��"O\Wd���?I��a{�ʕ\�+���ʴ	���'G�uoΒ�S~��<�+�zX+{�/0� 
2\�h\
�I? �܌�����﹛W�*p�p��I��Tc���yv��_����B4�Ի���*q�;�Ԑ�I��h~�w�Ģ��T�ƊH�i���Q�X�;��ut@읅�����^�x�1P�m�/OE�E����������i�WI��J �eh$�+0ܕ��5����Bv�F�A�Je=�����A�?֩��)
�h�I��)�dR�:��Qp�@zTυJ��^r���,Ȼ����'!Re�$�t�y$�L�C��<��[��:?��zT��p��L4D�i�>���jd���{+ B �HP6Q#Lo���c��1Y��N5��"�Yʌ��4�m؜1���/�����ޏ��[źy:�%���ar+v��ڌ��bm/;��Y��^����=��)s����,]'z��"
�?��~hxZX���d�D��S��}��3*���v�7��P=[B
&��hf쐰�Z.����"��Z�[�a���6���E$稈�1�"ٽ������K@C�)�k���dPkΈ�e娤D,��8I]�Ό'���s+a���^ŋҼ��.h�T��Lj>����
�(���/!`Q�[���=�|�}��g��X���O9�<�PH�ш0�h�J��Q��v��l�� �`!8��_N���n�k~�u9�s5�P%`v��G0W�M�m�:�'�6�_>�H"ϩ��Bs�� �5��k3��.��w�����0�a�\[�|/^:�.�U$B�6�d�;3��ha$@��r�J��|�l����g�4����JL�ߓ��q$S`P�)}�-��9_�~�Q?dt�`2�~H����P�M@?¼��@��H$m�]��T���\Q���!L�&C�>����w�u֤1C܌��b{ގ�����՗�[���2�9#��M���1�ԍL���Mtz�k2~�uc]�����'���Jlăz"����w|�_��w��1t3���$�F�i1b�\w� ��t����3���Hm����'O����ťBk�H|A\������Y`�!Y����WPD2����?����ЙfK2:�bdڷB
T��bԄ��s�/�����K�c]i����%o�*��6����Aa�v��Zv��ġ�!����z���Ў��s{hmw��t���;(Kk�4�}p�tns�쾚��C�Ñ���Bmm�R�eE�z�n�!9&�[] ��iPs����.��eD�B�}�]m���Gi٦*cXcm�ô�h��j@z������3�̛l��9\-|�@|��k�`��(?+Jr�=|&}�R;�K���7�_�W��5�}�vuo�W��Zؗ���'�L���X�1.5�A}h����EEo��[=�V,�������f�E��(����s6��9�r�-������r�"��H�k���xކ)�@�� ��'�?���ݥ�C�M�J"еcZxL#2E�^oR8]���� 2Uze8U=B�jkm�R��`�X� +K���������]gݮXpg�o��+��XA��\�������� χ�u0 �����vY]S魏�<������(�)BnD���zK��c�4�F�j��m�"	T$��zH�7���d<��N�%�p�Bs_i��Aκ�H���*(kq�!�3G��n�M�9�	����,h�����Y�,�|�	E��c�6�V鸥�O��Ǒi��B([�x�)Rfe[�
"UeS_����o7z뼦��,���x0�gKsE�Ō0��t�'�r��"r�x����j!�V$=ғ�@�R�|#�}�s�B��!7W�c�=8G�W�{][%W���_�8��X�d�n��E@�(�G���a6L�K�f����6�w��Kw��.�E���h!��Ԥ�J!�S�"���A&�����[��㷩������I��]Sb���q���xh.B��D��Ss"�+k�	���b�Rqi�V~@�uF�PR�X�'�7˚���#��+0Jt�D!�Ф-�Z�ʭ6D�u��ב����ZfPA[i5,�+ɸ�m��j<u��[�f0�����{�E{��?���rY��9��;*�:%ZUK�z�Ь�(�G��r���HAB#uDh3�8�E��˧��l}?�d̕���,|p39.�p(�>���pvjF���`�t�\P��#�Jw�2�P#(!S�/n���i%b�p}>�dS�ր�.�ǙBU+P՟����\�����3F�p�� ��Q�Z�)�Dh�4��ꃱ߹";,����bCu��g$��7�����DF��<�'��q�P\��?���y�ڼ�	���FL^������˲��>�>.Hf���0��4�R/6u�����=��7Y��D�P��?*?�$IƑ�l3 ���׏ݨ��F�zl�1 G��k���R�è#�k�&���	2&U�o-�G��$��"�߶3${�;�<f���n�A��D���dT����<ZP�G��p�>�'��A��=_|��⒫0�B��(�w;D�b�*e#����`.��ll��݂����RK�^�~��#����_�p���] ��a�霨f�"d��| ����Qٹ](��@R��ͼ�Ծ��	�Sܺ.�W�H�w�g��lz��h�h�K0XMϰ��6�'�{�#�o�"����N��ok����M'� ��kN"v�|`d��D�]n���AM��I���8F��|�r���7{"��Rg�_Nm�E�%a
�ey�v*\W��9��l�����}������f̩�����5}�K4LlM$��6���!X~w	��֙�l���F�n��ހbx�oh�,�*����냪�5�&]�F�C����.R-ok�C�/��3(�n��a���V��@N'�X'	j��u`?W���6�j_J��PS0�=��!o�����cA��/SM{���*Gp@�3U���&6�W4eA�Lo�E�t~c'з��<=h�䒭\�@���
%�^����Z�}�ڢ��'1�BC��ƃ�3� "�L=�C�ɣS�l�#�^>�n�."+�
��V�����}��C����Ď�w�$0�ɺ�M�)6��;�F��m���\�5���otක.�<��Pu�2�Z�x!� ���Z��nԖ�>@�z��מ+���v��;�"�'m�Y=��e�T_�b���ř	���܃h���Php�ǥO�P�0K8�M��)FT��P�&�D�[��������rGk����ga�j����3�`�F�P�3�F�I������k������֒����;r�M/NL*���x�R��%�"����2�a7�TG8�[�P��'�����շ�/kQ�\���dH�6-^�l����>��'��n������=D,��;�4|�(Q�H��Z�,�x�(�=f.�1u��k7�y�1tm.<��i��^T�U���� =@�Gy=�HK��a�٫o�{�?7�IR»���P4+�U/JAy%&x+]���#7�U�$���� 5Ӝ*p<=R�!�g�/�+B���=;�5(�`��·k�=#��� /�;D�7�8u5�8V�$C��/�UU3t�	䚀f�� ��I�j��A�Co��z�����tL��Kj��K][�z���x��k��m�NhwA6��\���~޶���M�oҏ�,~D��<�����s�)�����F�Rz��n!�:j�W!*�LpO��\Dm6S��XLK��VE��~���ۈ�3&C�L���CхAଫq&���9wd� ' �?�/)�;�:������t�0lA7T�����"�:
�?���7&y���*.���s[� X.9j�F8~@1�[D���}2���<J�b������S>�6	��|��#ȫzr�ث)�c!���X��Ԑ�vs��F4p�>�e�I�A�����"l͡�(6�ܕ,�ͮ�x�Nw��j���Ckѐ��xy�����/��@�I7�yu��W�g�1Fq��O7�<`�'��rϭq��9q��>7��'Z���LT!�1����n(CkMG�S�k��W�ROm\rɒ?�+{$������fECM"��X�$�x����Ɖ�衯N11�����0#=W���
�4Fs�A�N��P����"��(�4c�O܃,���z9 �s��q�S��}/�mQ����::���ե�i�-1�elԨ�Bn.MN(yc�����y�h�:P�%މ6�Trh���r�a��Z����N��\�9	W2Y�q�����)�z�r�Z�Ú��$,Q��,�W�Әۅ��\M�N�E]������]��]�������1`���T�}cG� ��qϔf5wT��x�S�ȐdOW���-Sak�I$�b�T�*{ (Hd��ol�/t�a�F4��q�X�H2c=ĝej��k�;GZ�y��̵%���X��[ػ�<�Z�5��˗;Z������V_}_����c�*���M7��ۢ����{����@#]Z�=���a���:[$�;��qD�ɞ]9�z(Wh�Zq�����̑Y�5��MQ�S�
S(��w��&~c��͙ݹ���R#�t�5{�����E���#�C����oUǁ�Z�3���� �S���¸�!΄+y�*���VU-`���vD1�>_�oLg3���'�O��٬&�7�i7�gb�,�v$և��c�~Vc��C��*�����tMȲ�T+�D$&߱��2���E��k���f���YСr���ت������ƶu��qf�Vߓ1�WC���}t����G�`yAW��H��������	O�m�-�^(7�	j}��N��G���#S��~#y�5��cQ������IYX�)o]?����KsՈR��Bv��ٟ�0�S@夣��J6�΢q�B{�N��b�B=��0D�ϴ^f�ne�H#�5Q�&�>~g�
������C����J*1�Fy́�.*�T��WH��%'��U��݇�x��ʶo�-A��l�pȥ���ߊ9�Jrn鰷��`�ϒkz&z�;n&&��I��\v-d<M����U)őVx�M3��lX���H��O!����i��bp���Vr�#��T�[䄑:�����ۓfO\:���7��~�N�nLu_���>��|���r����w��F�D�F1���	N����� �Z����b�� ��J���ӓp������ڕ<:źnkأ0OG^��ln��g�HvN�Q�����/5��6����)��tF�Nr��2!9�"������=�3:_��aO'y��Y��G�0�6���Odhg���,B^TJ��"��~�?��/r��M��R�NN��F�-�zh�(��P69N�O�'���Q���m �F�ߘ�\����s܀�Q�cg`M� ���b�O�\�����h>�n�����R����
�g�V��|�T�ج�~�F�g��4u�t�9��Z�s&4���|W�(��e8����7��M����� yʐ�2�x$.��C>�P�%� �E$��iH���g׍�\�'K�g�_�DU��Xm	�hw7�EC��!.�ާU�6�U��zwF��na4��&D�͐�Y���~��*F)e���Gº���Cn��޼ٝٮJ|{II�~��:�$[�p��'���c�0���2�Y\���}�4��Zj�ju%�h�@��k�~[q�T`	�Vh�ut����\�S�@��M�Y���H���`����k��x8�A�SN�+�i�z)��o�z{&���R���OS �a�A��[���;d�^ :Ɍ|�(?ө�0n�D��3DgF\���.��Rrv\z�fxsX�|0��S"�!�[���u�C0켃�j���T�8a�k��a�)My��?fzԛ)x���M[[Nl��,$0����%#�����:��S�N������{�F�F|k*hU����~r��)�y&JI�y3�1������^�;C��z�=���������0p����m����H$�U ���wOh-�SO09��7_p���9�ú�f��I�A�ٍEf��4"U��ak�wro�g9֕��c
�WkLXM,A���/��z߷�e*�Ɲ�@��Y��
eoݧ���S�����#��R��Fh�<3q���Xy����u]�vE�����M�gҢz�+N�G�"L0UX������Ky�j_��d\A����s��i���xh�զ�%gV��3�瀓{������r�|hw���j�J�3���C�yoX���j�����+D4����1$�-Y����<.��{9��a�O_�>�a�m�����G� GmՋ���C7.��F�	*x��|+�n�+S�����mk�|��+\�`�/׼R�_�^�����w6:Kx��]�q[�OTUf�*���R�x�I���d+;�Bߠ��ht����1� ��o�v.-�-��!���Q��Ew2�M�Z��1�"2����:!�e4⑿�C��	&��E{�!�v���(y��� ��@#d���0����81�iu���z�Ɍ��=iZ1�4�f���u�kY>�#�>�#�i���R���YTS88���~p��[��<Y�n%s�!Ӽ#�zӏ����-Ǭߖ�-�]��y~��D�KD�g��s:�\#��`4����h�t��k�X���?dO�8�±���60W��E�Mo�i�w�W��,h�
��?�-j�A?�����|�J��g�on�1/p/�~�6�l��U����v;�D�����C̆�	�.�5��t4�Ѷ�&�A�6Z���3^b�����r0ΐ�*֑h�dG�25n��|[���D| 
!���40��7'۔?^�5O4ƍ�������{.a��}N�L� ,TK���(�S�����XE��cJ�;!!YF�?���Mܹ��J:��f"S:�nYЧ�2�C�^L�u�g�G��C�o�A�9I$���K���.FW7�դm��9��O�PQ��D�R������B"��"��l �P��>���DF���Q�����wR�'�`�&M��h�4�+����G?���Zʉ@�]��6����������|�G�t�>��M�����8n��j�D�	�	���/��AkK�4����6�pt��<;i� �`~���4�w�������n$�lP�}�F@a��H�c��<M�$�V��9{��M��hh�-�ڮ3�++�.�������<b?{���V�����}�ʴ�uCfߵ��>�q�O@�j�Js�Z����Y޳u -��(�{KȞ�r+����Mc�I�+����\<͈L�H�
�	$�#�gs^�.�U�r��l?w(����,�y�]��ҩ�-WӔe��tN�6s;�i��9��qʯ�X�u>��e��~���Ȭ���T�?jN�O��#i��X�N7�2_ɿ�i�m>�M��'�wujjYm׊���EEd#�6��0����Ujˎ��<�
1^o~&e��`_���V��}'��O�@���l�~3⃟r��z*�O�«��C�W)u�o��a�*���W�����rO�7P�n��� Ҫqo��m��ԞvB��Dr2܃1�s`��iq���+�Z�9W�Eϻ�1�uJO���l7U��m�}�s�#J��ꮶqSL��.U�E%1�4 �-��Z�!p:����<�������ʖK�v���c%r���}���vUb:�k�"�y�*]�";ږJ�h�1��p�HY�t���&��Mʢ���J�L�v���b���2�i2O�zAD��"c�4���xn��8�y6=��B�X��TuD�̑�KA�C��vh&�jZu�ǋsi�i��7N���W�I����B��M����uՈ_�>$���T���7�z#�b����Iyz��+!�u�M!���0����J:d{,lwff�J��HU��<k��m�0N 0��4h�����+{ܝjw�������F�b��n�Ȋ9���G���� �������G��D�Wc6\Jh��1xy&�ܒk]-S�M��*��XΥ��
;�����'75#<C��c�G���\`�l�(z_S���F�u���l�$���j�]]�������f
�ڝ�u"M \`+��S��e�/��cY3��v̗xg~��Y��ޞ
� ����zˈʰnu�ɝ>�6$�vx���Z��i+�������s�jSs|	M����0{_��{aX��e��H�%��?�S{B@��v|?����<~��QG�x�O��,�yG>�{L���(%�ʊ���Mo���ŕ R�wS��TQh�$g�:��rL��u�yBTO���^^�_��w虻��f��͑���kFZ����;�V�{H��f�X�z��V��,��s�4��M��c�z �%�ZmW~4_zK7��#�Z�9��i�)@#������y8��UPY-r�oT��vmo������0�__��P\M|u)��/z&Ѿ�d�+l0 ��mMI<"AG"��H|��h}9<�	(6��A����������l^UE=�(�i���\��t>E"�}C�7��V}ܼ�L��U6���/?����%�Kn��00�;rF9�^*'Y�|�ԁȮ�GE�ِ�+�+�+;�T.	�U��kA8�Z�\jx���U?18�@4�*b�u�.��ĉ��_ ��F�w���ʀQ�O�:���+�#<|��ɷt�����l�5�A�,R	���c$��m#y�:�2p''�E��ע�Y)�ۉҦ1�� ����M	�	�nڑ��ߞ@��EI?����K�`����_y�%�D��m���e+:�S��n�u��q��{�΄�p��kb*��ύ*:Y
;�i��k`�I��f!%��������z+20�9i`�X�W
�E���n�얢y���%c�_	�ރ%�~������s���l��W�I.��,4+�4�!���<Yt��Y��8��*H����� ���ѭ��͡�ߏtvB$f�28����L'��M�-�.��]�+�0���=HEx(��]�+Z��)�i�,����.U�E�вA���"�T���vh�Ed_�pbC�/�lh%1��eNN��х�L��f.�r������l�;�:1�&қ��9w�
�H͎��s2��ATPc���"<C�h�vM;� &�̧���m��T)*y)I����h=`�o� Q^=-�D�`�mڣ�C��츷��o��yd%;�%���2�����/���7�Ɍ�D��<G�!a\�i�8�4�9��s��N�"��Wfh��5g���L��S��]F�������u��!�:SxZ���z�a��/Ú9]�Y9K�PEr��&\�1�����z�$_d�� ��{T�����d�rw���%�p���6F!/0����T���hm��Δ�]8*V��l� �w���XIrTQ0f��<<�\�v��}��{.u�D/�Zh��'��g��S�L�mS�+h��a��r�~���.8���9Tw�` ��1�꿸gq�Y���w	 #)5��F����G
�H��U����*�x�X�%��٦(�2@
˒��]��#���.fb�����+��܀��yٸ���[����[�?���a�t�����L���m	���ح�T'�b�:���7^̍��Ǖ\�W�ؓ��+b��=�iy�ݸٟS����`�|f���"���M�s�����g%O�2���*��&�r�\0|������2<���ߍ�j���������i�]����-+�l�B��s�L$Ӣ��3��/gU ���$���ǔ�ڇ���ô�v�����/ű�K��f�F](E E�*⊻[4�[��䍄X�ߑ-�F�f82x5�X���P��rz!�#%n�6�3{�Υ>��SU� v��|-U����q�x���X[� ��P솭�*�N�FdQ�tI�@���gL��О�p���
:'IU=ąLc�N��sw#ke�+�?H(}6��t��1�i@]�|���/y�%�w�y#�֦p�r�z��Y��e�ă���T���vѲ�hsjX���pF��\�pZD"�%0-�|\�#m2��<�e��<PA �#3�1�V��\�5���œt��#T���CH�s�a��&��"�_	��}&��(�:m��Mn6)T����:���h�cfq���I-Q8�a��	��$)���J���s+�$HG��B�x�Q�_(�\���޶mw7d7�Ϻl_�q����E��|{1����%�CGǛA~�LvY�I�!�;(����d��Rm(i�8��ਘA\Ր�c�-��T�諄�oa��b���a��9����q3A�P.��PC���P#��j�Q����G��B!��=(v:���[��6�FQ���Al(�z0�z�{~]2��z�{G���?/���jOb�XtOc�`k3	����L;S�ߢ#.Nwڀ>��"���fu�x�ʖW5����Ŝ�eB��:�i_���1V7�M��������PK��
��s�F�4�/�7Ù(t�d}`��.�u�$�A��G�@�g"�����xeӬ�*����Z��?t ��(Nv��Ԃx��X=���pf�m]��E]s�+4L|�}a��}��d	N��n�iqGC��Ka��G�5�V3����l'��\t�z�!Ty�x��a��x��ڢ'���Q�D���3W���54Y�b����Gx�ie����El���_ �� �W��l-x�)�i�[�$��\G�R-�*�F���9jP��x�Y�>�GgM�`=�t?z�c��i5:޷�U#�"W����S�B�o3�*��i����fn�bV�yMA3������/�|����	�)BcIM�f���7yCˤ=�,���;�c�xʳJ�}��Ѓ�������t~�;ǋ��m�d̫ ���=6�M߂n-X�|�"]_w�2��,��F]5ع:��˞&�났T��Gǧ_	Tw�5���=�x,���s�n����P�˖ޓ�O�;�?k+ Ů�H~G��厥�*��bq�[n�$�Y��P�?w�Ɇ2�}�*>�*����Ͷ[�9%�@2m9ހv1l'��b����C��3��P52�m�t�*�9)2�c9�c-���We{��b���pM�Z�׃H@���>Bߡ�1Ñ��tt@:^�x�0m��G�+}@�h=3�M��tծ^���f|*�J;�?�,kT�9	s��m�-3Ǒ~���^�b� *|�/B�K>S'��1�Ă�̽���~ƻ�Iu��[z<��g�Pf�F{'}��*��Υtl��H�Y;-;�N���5i�##��&�G�!�^&r�P$L�������u�K�)�,�@�Fc�$5����lm��DG))"M�'H����AK̢v�w�� �Z����7��~��|��J�?�b��^(A�ҵc�]�͂|/�Tr&�7�M��k�&kS��-HU1`��}ўٱ JU��r���~K��X�"�:�~�(�'�ǫ4Q*�v9��l3�u3ʁB��0�w^��)�U�N<Q��|W9F��d�
��T^���.�q�E��9`r�!_�$�І��{r��J�*ҩYM�&͏��N��qf�Ry��2p�mȨ���I'���	����ZR��^�:�+�'}�)o��6}��;>3�X'�;�����`s`�e��o�@�\LB��;:�0�M?l��x��dJ��Q�Lâo�b:�$��]���tii���z��kq)f�����zF|��q�-���x������[�Y'(����N$S���S�kĈeYeG%;��_����v�Q%�m��yM�cn��\�[��7k��R�i�����S� �0k�f�B��uN̓�=��9%g٫N�(�jy��J�F�~\�ڏ�������VƥJɛ�@�W�,�s���������q�T��y�
�����z��Ѹ����5:ok�%w$���*����,�U�1�<�Au����� ��Zݽ�����k4��K���M�b�Ad*3�9/��"t�a$ZxċQ�Q��Ƌ��Q�x1%FT���w��G�{B�'�`��.�d`3���	�G�� ��/ �t�6�?Y�@N���qO^{���f��f��q>�:P6~J�#�ˡ�0�SWI�f��#)e�7
��[��m0�;�$�<�u��W��Kf?{E,��n0%�`��0���C�������b������3���C���ǣ�@��^�L�+�ȱ`���꓈�Ƴ	j�׬r��0O I�M4�|rN}h[Dj�&T�ɠ�n����vK��m�3�$d���)�{a�֙���q�O�I7��-ӻ�A����^��ۋ/���ɝ��|�1��)���i�����
i�=��+P~�O���xw)��QrK��D�P4'��C�熄%~yY���U�&��L39͜$Fgn��9`�X�38��� ;��޵�m�
�`6/��.a�D�f@sޫ{�=�m�@�� =��RP��;>1���>��˭�*Z��}�&��K.�-���'�p��Y�^Q�[����/�Yɻ�d'��U�c�Ό�)Г#��F��]�6�N���맰�� ;3Kp�V���?w��)ɪ �Tp������d2?1����O��B���q�oUsk�q���B�-�R���wi)-�����<�˔��w�`n��s�5ȗ��^�ەW����ӌ��D#o�=`9eF�e��ՕМEٓl^�%ﻑЂq�$�*b��8��yT�!�D�F33�+ZLP���#�:� }���z��G_g��`TEA��a����0����:(0et��C�e�t��ĳ�|Q�V�²F(񫹆�TW�t:�I�:�)�F���X���l�Pb0]j@-KCG�r���fj��Z���Oz����:�v�8�킊��	9��02,�y[�=�&8
Yagl���طX\a�+�2a�SP\S�Etȃ�Gӑ�i ?y��_�\Ek�m&�w6�LnB�Xcl��:�:��*�yb�?�����BV�JeBmF�3��� Z5���C��hj�3~��{���AB5kg	}��K#�ܚ�"vp�=$NՁ-�'xs܄��E�l]�q�=H����ʝ7�SV� �$��r��	������ŉuh��g�R��Pv�btﱡ��@�(펀�	�U�v/)G��Ǉ}�-����]��_�\�$���F�~@N����@���kIƝT��~��g1��uIY����j~$��ӟk�pJu��S����v�ƾ��J@G?�u�<�7��{!�xFP���?S����X��'^�
�,#t8���x;�8�z��킱�qL!��:��v��t�7�s�zL��}�v�P���F�5��r̈́��܈�3Ü��1>�1D��N������KG2�3s�ݸe�c\pl����0'��J�7� o��Ry9��,�{l+�˙��ٔ���e���D�3�����ax�Լ�Յ��L���isd�$M��{�x����F���m-�8�O-Nc��!7$�c;�O,��uٺ(��
��o��V�`��k*��|�g ��!O�] m#Be��$��.'x*��,���{7�L_�+�t�X՜K�{���QaN�t�Gz����U�"sΥ��h��}���w+fy��n�E+VJ8q��9_��M�>˂kf0힀t�eP�$��x��>D2X�|:ԙ'>.Aӓ�b{��*�3��P$�@B�k��Ő<�,P�����)w��a�~��'ΨnJ�/ޢaMjh��D��R�����V��Wr��� @ԓڌ�b����>s]h,�leoDmSWC�x&<��:����3���F��q所oa�d�Ӛ�0�8�H�Li��J�f��<�*�h筥Sj.���E�n}�J�e�dF�YLf�bR��:��"%TXb{P<&���3�*�/��F�����(:a�ױ&��w���ֲu��@�,��`S�N�S��=_��Z�~{/G`���`|�~bߨp�QTO��h�O�uL��2Y��f3��(�ߒW�����ڸ���NT�{�oN���a�����B�!	K 3Vg*���b����׵_�\Ϙ�N����Ң��IHwٰ����ͱ�G� ��	�z~�ݝ7�0�Fw��-�"�w`���O�&�ZIO�78�~�y*����. ��?�ة��k�OƬ�i0�b�/ڼ���,x��{��6���$����9����p)��r7d�����c��tk�^~�y�b���RJ�)��S�ޘ���u����!&%^�[C�|(���P�����s�;�@y_[��[�_ի���0�^ҡ&�z���BiS)�.L�ȯ
�	����,�G�h�<�y����-�.-�XJ��W*��SS&:�iP������X�U�@�`'XY�U�m�(��@�-,��1EE�(Q�!��bn�N���*^�13����:	������P��#e�(
'�a��~�]�i�W�[�&�1�\.ڕ�]��\]-�� �����y}z1�7ظ�Db16��$�#����UB�T'��!I4 3��r��+e�`f��N�N�y��
�����f�M�"����-lV���ߪ���ksH圓c��w��7u� eX�a���R�'~���FC���<���nj-)E�Y`Ɛ�f��\d�C�Q��1�p0�	�d���#�:�`ڶ#����ݼ�te0.�������a�
uI���<�z���e� Y�&�H����g�vrʣ]�&ޟ��s��Mr|Wc_���4�oF��t�Kd�b��-/_񅛋��CD��7���Zq�4��6�dhe|?`-�Y�,�1��
�i�V�rVTq3���O�Q�^|rqI��-�\T�^0Jձ��r-$�|�Vg�$kw�#��TAt�P,fm�����ч�nv>6��9�;d��_���R0J}˅���*6=o�7�rː�;x�9��X e>9^e5v�$���	��G�]�;|�%�k�s�1T_�m�`�1<��K��X��׌}S��9	�p������m�A�bS�����`��+�	�#8�����7m�@��@`l���HMWAm�;����Іnŭi0k3K���&F�x�H&_.����O8g�\Ere�M#�Q�����6 �3�ν��u�����͈NB��tA�p���M�*��b���~��f6��a�,`�C�9Z�+`�/��{`u�S'�Ĳ�am����{s�V­��+����{��̢=�[l1Е�K���pU�py��у��h���u`JgfD�T2B �YM.c�Rʹ�8��_�k9���{D��!�/���G��z�C�-�mA� KN�_;'���J�c1���;tJ���opG��bFU���!I�ףK0��%��#I���������@̻�����>�pum[/��<Ց<�w8 ���b�e��D2P�cU��Y��eK��/+Թ�(��;�t��̓B�O�VZU-]�=�����OG�g��	=�x'B�	~��4on�n�<�_Cx]\U8V�
��1r�YR��w�������_r���C�l��1+���aJtQ;L����5Lz�Z��0�����HU��
���V�u�1vt_��<]ݴGX�^9�^�(�_4pY���<�U\c$f��|��M���d����U��Q��}�r���tÇ�jV�*�Zq��9a&]�ȑh!Ѧ[;�QC�X= VV�7�'����ǅ����(��S��]ndcw�D5�-zVp��J�t��@o+͔o]�q����,��7�$C��,��4��	Ud�0�J�H���e�J�y���Z�w�r���fȊ;D(�P3�17/����o1�s� �;�zwR��n ��<3�8��ql9Ps�c��B&�˂��Dv\)��2� �n�ޤ2LCAݔT�[���{�a��j�j�,���<U�ی���4��^�Zi9 بA�FFGڄ�UϹ^����Cz}¸�Ǳu�yg�$(Ƶ*`�_��؇ ����$x\8?tx�8��E�^T��M`N܌x���}0����x]Y��g��8���V�����4��	v�^ὒ�k���~�m�� f��TT�{���Z<)T�|��߆���g���*Y`�&��lЗ�\�A���u��NS�Zl@[����IϢ�������\0�siۮ�d������[׺X^Q㇒��[��HKd�L/��H�s�e^!�
�@�9�����Li��Q����� 2o�t`�Htm�l��[�O�^"KQ�pUA*ߵd^.�:�8z7xX�*@|�����'&L�_��">�����JG�;��LE�3ߺ�0������"�Z`��(�2`��TrI"���"&k1_&:��љZ���݇�n�nL]��a0{�l%�f�Wgw��;S��*��I}�x�؄i�{EQ�t�����׃�'�h��wdH���I�N(�ĩm�)^aL7V�(U}iA[X��8��#�L�[��Qm�_~ب���3��e�g�5�w����Ay`���p��?J<��u�<��#�l��� jyK4^v_ˋZ�{k]�O��=~��nx:�k}خ0t���ڀ�[�_$	?\$M�N8�gU�P}�a����6F.F���N�ø?��������^����W���� k��p_�r��o$�+�)1:,�Kg/��ՋR�{��-�����\풵N�-��o�JI��9���2(��R�[�q��?��P���d�c�&狷��y]4/��0���V>O찉���oڠ���3��Ǽ�M�ן�]��=�1ȘΪ`pr񤺥�A_V����v�s��sL3\�_���E��wց�GFE�=~��RUu�����5��8����ga?���{	��(�j{=�����*�v:����y� ���H�mJ���o�I\���O8�k�������MP�3�9O,����:�j����7.!���%�L�Rb����6�ASd"I�L[j�2𗾡g~�1S;�£��p�Ϋ�N|z"��h�nMe����(L�Џ#�����I��i������_�����X�����jK�۰p+<qjt���]������4��@A����NWUp�����Т���pge���i7��wy0+��� ��Q��X9��?B;;Ȣ�k������ �Z;��	�Ŗ��r������g�B	g����p�+X�ɩL��Ns�|uhd��I�>�(�o�籱nVM]'�p��f���#��^ꃣ�B��A8Ϛ:n��/{X#V�
����FI�9f��Sb�� ����͖շN���H<#�yO�]j�H&[熞�m�+�N4[O*7�Ѣ����YM`=�q��y �3K =�QK�	�v�8��� \o-�r��%o*��+����R��Ƹ%��x��]�Y	��^�5����.~@��>��|Q��:W���<�?��̠�-}^�v[q��*��$�?�M�6���`��j�p��-O�Ɉ��K���1w�=c� P�ʓU�̧�VH2��&�s��ԚD����"�ȵp�rm��B�<���v�@�bxrYk>�'���Q��T(�ѭ�-%4k/5���Vި�X@ �����=���N@��g��ZX�΋f	Q�&b�-�"�P��>�V�J��{Z���3�cĜ�3q�T{�߈]�+fя���'��V뷿�{r�ˎ��̸��}JZ�("��4K7�8��'�͛�>_c6�K���|kY����L���_6�vaݻR����ʙsX�Q�k��Ʊ�%�_��4V��N̼�a������'�V��Sve�]����y�`�Y~���6y[8������"�P��͢E E��ĸ�5�x�p!��k����}rN�^��O�f�� h�U��*��S��c�A|)� �	Q���o)D|@��<5�YQ�6$�}U�R�� �ע�@㐞��礳Q��*Ҹ�4tO{�DS���5��I�~F�ϼv.��!�:o�G��g!�v�낈�9ng��Ԧ|�eA�k�8�!�<!ie,i�:|�e}����i�����C�(Bf���{��4�Bۑ��#of\��^F��ӐR��[j��>�`�髱�����P���j��;�%�~��H��Ыe�+;�
�5���P���Q��`KLq܋���ř�9,�T��2QP?R��W1��4%�\���D�\��)	���N�܉���ڗ�ymH��I��8,ˋ�����J|D��b!�.ma%����翃�W�q�����cz�N���2}�!�gqKǑΡ�p�!pF�(�N����u����A�$�V�Ҧ�ϟ��;=\����>��q�C�����ZOu8]u���7�e�n��[,��SCY&��M�5a,�q\+�I��b����Mw���2|t7x�u�����k"K�_t-I�؎M@���1�=�s����Y�L0�)�P�Zd��y��3��6��}]--�J{;�R��ڿQ�b��"t��<ܠ|�
w15.�0NZU��*���W*���k��L�C+���VCVv�B< (�~\%�v�W���Q~$P�8��P�W�g�k���;��YK2f�p�J�8��%LH���ll��&s�z�Q|��$�K�<�+y	#�/?� ���?�bY���R�$dC�5'0j����&y$肏�\��L��z@2���Gx�3�>���D!7���Y�f<����lPF-��ąWЮ�����Aatؾ���W���E>�sz��6�yc%Z���{٣��j�h����7;��#(���.ݱ?�qnKX�]�f��+}���徾�vL�%�Ҥ�s/L�"��9�V��!��x~�_y�h��U}���D�+��v&}&�p�3��}wK�h�-�z��P��0WA���m��k9=���<%�֙�[����M����n5��Ș��g�w�'�y~ʷ�nZ�f���7�����q�Xg���7/��ߊ�bgA����S|M;�EKu�����xg�#��ĳXW]���f� G,p" �c[�F+�MQ-���\�#��}(`����ܵ��g����a7��t�ȏ�hI{����O�	�ʦ���Sʙ5������:II��1�f4-� ��jҠLň�X��	���^�4)�a���z����?�d���������aނԊ˷$��hE��K�~���/�d���m�tw���	�!$�4\b�;O�i$m�������T�R���!zB��:3�ڔ
�������a��B���bX�ǣ�}Qt.Ǹ�_�ΨD��_��q�P��Ƹ��!�a6�f�)�Ad֏˳M�l��2���؝{���f��,]O*�����fl+��I��R�e�#���	���C6J>c�y��3P�-5+U�\�����s\�V~V��^�k�^�20�U�<�Ȼ��[���xZ����G��{q���$��k��8	���
g(��4祛‑�j�rȸ�a�
ЎM]D���,@����.ګ�2��曥߫ٙz4�9˗B6W�?]�4c�淶9�,pd��_,3�0���e�W�wOD��i���)�Y{h5������;Ų�~����˸U
#?�W�7}�ɥz�B�ػV�g��n:Pء:^Pه��

P����e� di�;�7�(bH��C��G�r����L�E]׳Ժ\g�{ή��m납�p�U3B
UE��p���"pl��� �i/��K&���e��z��z,�=#�	� ~���m���;Nוp�V0*�'���~��ݫ��vP��BCyad��y����$Y�-8���e+a�c#�ea��uUy��m";�Oȧ�үXt�eY������+�\Z���R-9ǩ��A=����p�eLvB��i���i������s+�@�m��u]�0�����ԩ�<�#�r��Yc_H�TY�!��^v+��3>��s+s��K�v�}�_X1{%��eKj*F�=�՜��x�H&��CT�v�,a؁%�o�!d�!R	A�_�৺6����>���2U[ddC�l�^��w�řZ���j�E4`��$�=�H�w��5L���2�
8Ho"�6�|f��4�ޫ������q���9y6=E�V�����A�dyC��~}7�֎���������{�|��N����tL��9�Y[nq��V�+td0~ؘC���;M��l�;�e
`(5�}y�p����� �!A��r%"R겼��!�8?�ؚ��D�ę�4�����Dlt�4J�lпH��l-���J!3����N�+]�����?J؊��̋m �E��j���V�|�0�/�&Ü���R���!m��x'�F�Z���d�lb��\�#�i����9J^��3�v��E|/:�R@�L�oC}�<M\/��WN9;��L��0�=�A�3/��t����AH_��O���ԣR���SUM�+1٫��=Vn�\�"}��t�y4P<���F��g)�	xZz��K&"cR��Y���ߐ�˟y̴ic=�hD��$c$q�/���sg�?^�V�=��aL�P�<i_,5���9�L�ėr���b���Q++�#<2��m}�wz䖤M�isIY���X�Dh:�B55��dC��t���[M����f�.�R��0�n�_��XRPn׬��x��a^�"�\�� �HK8������o�N��_z$h���0.��s�7��<AL�`(e���c�,���5R)t���3d'�/��T��x�_�~��OL�]u3Y�?�b�̹t�ϖ<������b\!�g0}U��c��o(��ۅ@�Ji�w�,���`�	T�lK��w�gDuB���W��?{5O�̧߇Ve�C(74�C͌������w^F�W#Sg�Te������5�Փ4�ɘz�4���6'���j�:�=�|y���~VKvfD�az�I�/�ABoX�=G�d>�r�V�	,�(��4'��k�	��zBo�@R��.�B{O�0��#�x`��nMO�������״-��Ǐ5�����������#f@}_-������2J�c� :�$&ߔ-G�j�H~F�օ�´�4���*ϱzbV��G�m�>�X���1��L�Y|��d���cl�+��FHQ�]X�P �_!��u|��9�����K܆I�V�yERC��=W�7oR>��{oM��ќBn�F��*�Z܆�64������N����W�&�^a�^�,�7���-�J�x�"u��-9�@e������Q�h�7$J�����t��Jsۛ�_�dND�,"I �HX�`���E����b>s���"K�4�~z���^� U`L�$d��9�@��Mg���d�lC��7en�N��N� &]��(<���V��r�e��}�-�u2�U��Q�,��O�(�@�&�����& �2��Q�����O���M<��j�l�tP S]Z2������[p�.E)�Xk���7s8h�*���]G-m�Ge캪���*�g�M�Z܎�ӝ�F�d��<�eٷ∭�J�L�\����rz@�#�Y��X��Er���k�9k6}ӎG���-�Z�\�sB�{�N��B3(��q�.I��y\�c��M�	����{���\�܍�Y��'N[�p��A��Fø�-��TyɮHO��h�O�f<N�����#'J�ಲ��lSl5�M�}����Դ���͌�X΄�_���d�~��	����z6F�J8���ͫ�j���D0ݒO<F��IYS��ߍ^/��r�s}Z��S���G*�'� ��t�s�n���ă!�+Ecqu��_&�N�:l�K�r4�Qt락��ŷ4[���.
C�UF�5R;������b;��V�Р����)5hn���O,�#�ei��a�X\�¡O��IZ���~k��#�=2�`H���:�0+V3�Tt�B�m�$Cq.h�e�]MO�X W����-L;>;��E���rm=��G�Z���5�a��؏0�b��'���2"�/1/�[x�\߲K������4�oI�4.�0�L$B����]�2���_&A�х���ܷ9�X�A[����_��L�Z��; ��v�9`�t��B�|��?E�B,S^���ˬ}3�AL�a�xK�6(IO,'��ט�ܔ��� V�/�奼���U�,��|D8��~eK�	�v vd��1�8�����%j�J����.�1�SK�X�Κ����VRf�'��fBΌ��ws%-�q҆h9�t,:Gn>�L9d�֩�G&��<E���p+����$6ǷM�����p�ǯ�[�#\��oy}��+���U�]�^�!�Y(L�>�Zf-A>�ѝ� ~���c\jHJw�e�sM�qB��)�B[��V�� `�����c����徯M��Y�>�
�܆D<o�>�����
c�P��K�ҷ��3Zu9>+��Az���F�D��H�}���8Q}A�57#����B����������8�m���A늎w��P<�l!-�Ӗ h+Z{��a_��K}-SO g$b�P�@<���<�:y�8�a�QP������-��*́.QV�﷍H�8�!�mk#M�Vf�x��}��!z��\�\?}���4L�}�F'��xK�/]_�|�w�Ԣ�}�h��$І�����@�O7�nC��^��*J��+�޹�f� ���4�"���4����+���WB���q�V�:m[݉�c��c̭��L�h�dU`}+fbE� \z�MF�7��6=E(��=a�[������|���
�-�h�e^��〥Q6�@eI���1��=�?5�|@�G�*kbҮ�1�-!�ꪣ�d�L �4y��Aӵo�&���xB�QO��Ë�3�F�aH1А{��<#���1��
N�j���.wZ��e9|>�p�t�o�;/�7\Qwy�an ��"bp�������bl	�M��o<���DX��WL��}V�����챑�,ED���m}�H��ښ>S������A����U[�������2W�$6�ul���3�	�����Ӥ�x���2C>7J:�;��DN��؇3I	�t��� BR�� /��5��>�sd\���s�@k��}�Aj?�i��nj�g�i͔�U5USYRm�5j�Y����R "5��Ŗ<ɗ���1��9T6��:�.��\��5t6��W��@�7�>Lo|| ��PP*t�Ӭ[$�1�䜮�3�,�5a� Z��Ml��B�*m-�29iԕ�����}�X��;Y�Y<�qܙ08�	''v�M�4U�
�s�S�Nl�*�I�n޽�5M'�1�ڱ嶘y��,�6L1��+���5p�3X��+�7����hSz�/�z6�wI��'�[�k��ԗOg���y�� ���ڸ���@3q�~�/�{�Yy{u�n��iu,�=�m�I��lj�I����m��N>�B�s���c���	&��_^�ߊf̎'vR�����ìdrhC�r/�rz*<QOb�U�e��%�P*k��`�i.?Fw]��4���d[��{�i�M�.�3�]�����g����դ%繪`Y񭧛[�4g�p`����f/fچ_��qwp��`�r7�
��|�-KĘO]�r�����A���\��By�����(U��C���r9D3�'n����T���A��v�R~:yٶ�p���l5�V?q.F$ ;%�oEgxA
���&��׎��l��j���`�������hS�se�o�����L�l��#���j�02�'�!�4c�Q�4��_�'�(�4��M�>�%��NׅΖjh���}T̾+<��$KY��l�7*@̥���-�q:�3*-%��@$�qJ꾶Խ�$$��ȣ(���b^AC���_sr�[���!���I�?�&� ��(�tzN3h�H
���w����|s2,w�YӋ!�s����]0��q����s�s Ծ�𯍄:�I���DOx3�G&��!ғ�r�q�a�W~{96\��m����i^D�DP&'��p|��9������d��81θc�~��i��J|1�@��q���WL��^���+����;s�f��Yz�;X'��P4"����[�6��hX	��F�.<T�Q��p!�gVR��#]��G�����N5��rO�)�`|�fo�k.�g�KSX	����m"B��'�3��gk�I��
�oXN)~��Y
P�{&K�5��D������mp����\�D�,�7�wX����Z�=����M�|��@˭��,�*����U�'�**��:�}��dΩm��>\��s�k�0\ӏ'���է���ع��<�Q�˪�S�?�9c��N�nJ?�HB�G����0���kTÌ�On���gy�R[+�7��w5��n�Ǚ��h����K&F}7�?�~�١xD�E��,1<��/Q�YIP�>2X|���ώ�Q?�Xb^�W"�\�\�=�c{�r�����Ђ�d˼Ak����2�?8�9��߯`Qp*-l"�<0r��k���Zq�Jw�GF}}��+Q[�^�>�X#RH�dF�F���xl���P�ׄ��Ň�G�`Z��`S�V��,�n�­9
���O�5I�bح<9�5�{l}7�U8��q���j�iK���L+���{+�1�q�G��!r�����&�'���/�hK��/�EQ>	�k���ɞMу���v��)����dG.�'��'��-6GwH!Y�z�L i�;��5��,���MC�eȌCt�kk�G�� ���_�]��K��]�S�@��:ou&\d���ߵY�%CŰ���4��'�%���������&nE��A0:"�3�y_�zp0m�1��ى^�[�l�bZ���ܾp�(W �h�9��y�u��N�7!M/��K��0���ӆ�ˎ(P�z�>T��� �JD�UT�.��ۆ��&iV��`gb���1��G+0�ՆEu�M1c���Xٝv	D����v#�4�:�兦-FC� E*����e�ho�|��^���� c`"`��Z8
�t��S�����D���VcC[:7���Uvx�[�F6#��#��"
_^����F��4V�`Q�=�M��X��N�m	���|oG}��B�p���WE��쿨M���)j/|QW�������e�9V��(b@�P���Ӷ*a �i�$��ǂqN Y���v���^�}��@f8)��J��C&��T��[�|�B����J�̭��Bf"�n�m�(���Zͺg}0�W0���:����d��X�	��~MT��ڲ�5��i��c�	�e*~WI�CZ6���Gi(�g?]6b@E��������Y�e?xRw1HH#��Wy�H�!<qP�b�jW��)��i�=�x�mX*Y�vD�
��>�14^L� ���o�Jes��Qp�N��*"��O7�cՙ+�Ϣ��#Kƨ%���H���6�>�0�%F����ֻc�(N������ ���(�s}���i�@Z��v������4n������_�F�|��6�p����+��ۖL�aToKŉ�iz_^�0��%���:��Mn��֔2:l�Kn�A�:R��@����"��R(
v�9�Z"���i�2�a�Q��xK�@H�̅R�}y�����텋�(J�����D�P��L&�K(���[^ �Z)����¤*��'_&�F^9̞pi`��ϣ�Rǎ�-w@ ����XSQ�����&Vv�5��->0�|��@\ep�&�Ϧ0�)!�Z���F{x���O>M|�i1��2������T��
��X[���za��;��0[ v�姰{�%�o�U�O����Z@�m��u���a\� �V��5x�s�Ƿ�ͅ�g��mJ�~M��	�Eq�f3�O��?��v2*��YfO�=ސaAH����(�L4��< ��*+�7n+|[0Os��5.�5p�{�Ym?��?s�l��z�a,qc��48͈��h�M5��M,�AL�A]>܅�"d��P܎��ץ^�0C��C��tX-�:L��&]���*w�uE�Q�i���(G�� �}�Y>_�A���V��ԶlQ��r�̲wZ��X\!��!��6�nTx|������-S��V�����1�Є�5��	�p��J?E��bR��2�����%�E5����Z�yZ)�<�b�)����z�!i�#����5OT�����OM���Aܻػ� %��z��T�sӠ^�;��)L��̍�X�̩����:�=���(Z�>��6F�=J��h�O�I����4\!J��ƃv�خEH��;s~HD���ky�]��ς�I:I>��m�f����}/\�mE5+��f�9�I�Y����Ŵ�O��g�����T1ڈ�\��{V��K˳�a�x�9,�J졧ѽ��^�E�B�F�Y�}�ب�o׌'U��l�V� (�c�������z����t�������Q�!m��l�tx��'�C�'c��!����O")��1Ss���n��3��B�r���UbdHQ�Tw���*Z�mcJaa��%��3h=3�W~��(^���כS�x�������
��N^6�p�
7n
��7_��54Y�;�c���7��bܸw~[[�t�7&Nܥ��
*s;G>�f�R_i�C?,P���j�?`SE���Pԣ��h��?���p�\��$��t>�J^8=&ۖ�o�hr��D�k�G�ᙺ41�|���2�VY'.��4���.���U�v��x�Y5ȿ[f�Lc8Nb�f����X��z�V�2��D#�������Pm%����a��6��
tkQ���o��s8(Y���V��S��.��$��1�-�����x�CR$	)

T`�͆����ϓM��ͼ:��ǫ���A�C�+K��F��n��9�;��.FL1L� ��Xؾ[}������
ȥ��Z��9�%�0��|��r�s)�>*k���H ��p�p�_����s��W�$��1o��0��c�lG��#_�8�B��QŐ��pо�7-_uU��XI��}tH�� !	�����:�oM:��K��M�ttn��'e�^{O���a��0+�aJش�B1a���Q��(�Oe*���o-l�[�o���zM��������P�K�j�����M�Ē:�+���jR����8��Ϗ��ӵj����c�T�b���`/ ����H�{�M��$a3�D�R��)+��͹���9C05nG�Zr���ܿ����⡭N��5y��V<O��~'�ХR6��UowuE�fr �:xH��1�!e}x��ׅ��%p��ؘ��c0�B��3\a��OA���ln���W��R�H�b�g�9HsǮ�I�����o-[ŃP3+ݱ����S�('���?ZP�������ܟN"b�0At���!0�*�č�\`�D���`�~&������!�B��F�i���¹I��:�e�³����D0�_�8{D.�X�o�Ҕ�����;*�mp��g�%��Q������E��D���� ��ࠊ�/�eͿ���ə��6� 1ئ�����ф��RG�8�¥R�Lyۗ�,#)Fzх��|��.e.�kjy�~,'�K!E��.�:=���ဲ�s� @.=�����=�4E�S��!��[�w�b"r�V�흾-]jO|�Tg�����˳lyL;�Z��'ǋ�Nm��o�Uʝ�K��.Zv���x��~��&�*ƅ���	T,\���(���%��7 �s��w����@A��7�,P�~��Uq0�U/"Zw>>��8c�d �]4��\N�ЙM�2�o��DI`G�M�e�M_��}:!�`x���� ]�ދ�e�߭Ғ��=5���3���ˌ��B �R�&�4��3�^�=��ӱ�N�������n��[ӏfV�Ik����g=��ri�������{�A�c�ֳ�wJN敚M�!�)�(�	8��ʙ1 I�U��o��@��D���#;DJ31��G,�E��ƀ��%_6L�n��`֫���\�����I�j�V7��LsR|����6m��}�R�	�UWQ����N�A�P��4 �8$9��^���t#����1ª5�6����i��X��7�����F�O���� �IP��uY2�6Q��d-T�(9�:#�N��J'Q)������wR�v���H�_33~�im��Ӆs�pp���ըG3w�v��b�e6l�ꔂII#����nk���|q;J�zOV��bWH�J�W��yo��)�nb֏��^}9!U�k'�)+&S~�I�c�9�VM�P���ƈ�qZZ�G�Gc�L�_��o3&1f�<�cv8�2#p��[|A���Z)2M���k��N��N�ﴧi�R�n�o'����R�۳�Ԛ��C�	ar�v �|S��aQՁ[=��gf��Y������s%�""r���m[������;Y�~��ˌ�4�Dk��۷�� ��/G�ֈ[��e�"ÚƯ�	�#e���0y��SQ��:Zĺ�����@���خ���1�ν'j��0Ţ�M&��^PA	E���2�p�X��	�~TP>f����$��"�����X�GP�X��e�K}����G	N��pƵ{
��5*YtX��Չ���$X=ý�M�|���3O�̯����r�A��*�`�����э�D8$�	��_e���%yS�Wܞa�ל���)|"f�a7t0����{��~"�Vs,{�J]��Y���(@���i�I{��g���6=ru��8�8�U8��0���'v�J���A�@�����|Mm�l$�9S4Fg��I��vxq�ޖ����V,�L��仙��u���;~����;�'�|Ы?��K��/����Hj��<g��r�-�A�,�&U �k�!����Tt�w3�HV�\|W���c�??��~�o��iH$J�H5R�
��3"d0D�����ȡ��.�6�MýQ_��U�=�m?�%�˛�N��ȣ�hn���W�����&�;6Zbʸ��!�/�G][�-$䭽��Mgc�f?2��
�qM;����
T5���6r6l�)9��r}�6�Ѫ�św�<�O~<�'�xJ��py�CsE4�H��
��bހ0y�.v/�}�nR�~�?,��G���ˏ�otƼ;2�o���