��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_K[��X���*���[����%��d�ۯ����j��� j?ϱ����z2�3�Ұ��j��#��Z��H=�dEMFf ��4G�n t���*���H���S��Й`Ol��C��m*�R��L��i�^fa��=����y� 6�w�a�
WY�j�{<�#r�w�~]��4T�C	�Q����u�(�^��� 5ѡ^��蠎�nx��v-�a��k��bZż1!lY�K:3�uHd;�����5+���^0,T���mD����7��Ocv��A�|Am��z��i�\a� *�),������0�����p��N6f;U���Ev=H X������#^M��;��P������י�s��!��"gK�2���^;ݺ������cb]([<��� F���6.iƸ�:��@P�n�)Z���U�Ju�k]:|�e�^Z¨ھ�{7&e�@�C˺�ѥ�Y��_C*֌=ɢY`��e�we͚�R�}ѽ���
BN1�����,ۃ���<�Fk#<v�����A�r�vc'f��YT W����H^�7��oJa��a��y������GG����X�ʉm�,t.p���I��� S���Z����3�r���b�M�����9�J��iU�\Z��;���7
谦G���Đ�-��%S�x��c"@+��310'�����g�t�4	�J$�C�N���p5�9S��!�*|=��&YU\/�A�&m﯒dc[*M���$i� Z+̻��7�<����#����iԲȍ5ڮ�)ac�n���J�f��I����O.=�Z�L�L"�g����q6?��aׁ5��p+&�?�pOJ<���4����Ee��r<�����l�����6�B�sMb����U\�E����25H�ٛ(��d��P�z�BS,v�(ҧ[���U��	�f�B�,"�-���h��w�'	5E�"�p��1�|]n��E�7�	\d�N�V�L�JAN3w,�<|��$��t�����&��8i(.��3����Ħ�t�j�*d+�V9�7j��SG��y��m+�Mj�^.��nG�3~e/�
�˞
��\���e�r�ϥ1�z5�f[�M��Jr�pͻ����
����h�Ʀ���u>�aI����(O�y��۬P�"@�6s,zYy��\P�2X�S��.Q��d,G��ꮂ�^/(�'䁶[>&\m�hJ!�O�^��(��N��NI:��)�ƌ�a	A�m�u5XBzi�9\�<���7�v��I ����A���zO��(Dz3P�C3�_s˗n�ZLj����*���A���5�y����7�ذ�����E��E1��'�9�_�G憥�����q����lĐ���-��L�/��aE�M��)}�j�~Qz��fNò.���I1&��b�-�l�TpY��F��9����źqv"�n>�� �]�fg|�,��#r������0��6Oq�k���/�LmJ@4�����`�FM�m ?�e$?C؟�bĞh�V\�Z�v�'���vv��Z��H\x�xv�#�]�Zk����ZFє?�:���(�bvBܣY-
b�g�Q�C�5��B v<':�Prԇ�c��h��Z�=��15�`���a�mx��6�T�H�,j�xoA�t�}�G?1��ܪ'��ۢ�J.�pz�EAe������O๽�9���|<���' Z��N�+�R�=�x��\�.��x���m�wf�6�'���vl߿���^�#��>NH*n���j�1ߦ3�����>�U��G�'�7�_U6��'��!o����*�S�� xB�jʨr5�G���dA���@;��F'+��"��>��E�Z_g@���5ٗJi�|rpoJR��g�����K������i��Wꠅ���^��~2=�%�벢Vܻ�	�b���D�m���y�*�D��Y���$�ripm��O�s;w'���.Jq�;-�Ӻ����Hs]�}��ݼ��1��i�1l�������X^A�L�7橭@�������_D�m�1�S#���6.Z󾅊�0C.���&L�����&q��a<�e^�ڲI_z�I����I��*,�2xy!�˔9b��&jԑ�р��%��Z*���磗1p`��������N��#���! ��Ʒ�����	���j���x�U-�u�>��t"m��0�~4퐍��hr��f����flV'��w��S�j�i�-8A��s��N�c�y�~�D!Y�����䛁��@��|�F�s��~ub׬W���q��7��,�'�Z`���ؗ(������V�;߸�ZZ��A��M�Z)s���K.�'���(����� �?��F;���dmU����K�PT,@���?��Qa�`>�0�cp
KKV/�߲Ʊ(�6q�Q��@`ewJ2	��X+M�SI+�ZGa�s�ت�"a����$�@�k� �����o�b�x�L��b��5�0G$�� k�唔�`�u��w�[��cP8ۡ.L�we*[���Jy&���YP�ٞ�~���p0��ؿ�̔~,�,�4b^�6&�QD)~J:9�
2W�}\k�Ԕ�2I�)6+�Ɉ�M�z{�4e�#�kQ���^�Z�1���E��.)��D��[��r�
x5��c�E����2��j�-Cu�\�['լ��#�	�]|'*3���̣}OӋ���c����$���$�q܀�!~�}  �We;ѱN�u�rX���":.�T��p�'z���K��Q/�@a,�ԁ3-O�����V%�$�,~�oŪ6�CM�"��/AQo÷�K<i�.�G�g	��Gt!m�X��`��:��X.��Z�%�Ow?�jn�u�����g����#:p<�%����ث��O�{9���3-�Z��2??�x5��K�6(��O��3~�Wzm3䱌s�N2��l�n���D�V���C�r!��Ŝ2)��˦�*1� ���񅖙��O9��C�.D�/��ױΞw�0���H�ةM�4�����Y���=�Zڿ_���1a��� �%�����ܐ�JTބ��n�tfg���oS�:K��K���`{s�dt���y~��'e�P��@������ɓ��-*kЖ���[�C�4PRׄD'x�8�S�<R��Oc�U��m�hzw�s*��`��F����2�)fD�}`ģL_ݙ<�9]Y�������F�4\G��hsԦ%Fŀ[tΘv�X�K��k�g�
x�lJBU������,��`.|���ɦc��ݘ=
���+�� ��t�:�Z�+���Q/'oQ$�`�P�=�*(��k���0�H-�nvo\ʒ����{2�Ȼ�6H�p��k��q��fb�k�R)�����}����A&oJ�V��=��Hf�}���82��R��s�2����J��h��(ٕ_,�O�?��-�����-sb��-�z;�����U˱����&�	72pu�G�ns������]K��(c�ӝ�[�|k"��e���o�C�B��ɔ�\�Af������y�Z���� ����\�D'��K8�Fz��>�O��tT�Y Ѭ�>��J�{��u�ۙ�E!uYT�ut�\���S��#�;�JEb��a�n&�]�:R��c<J�����#_�b�<�*�6�̥je��,��]*����A_�D�w�W�:g=l����n�R�r�G�/+�Tc�B(�w���E_|+��@�>i�k�h`j	=����&��Zy\��B������Q��k��Zx��#�d�5p��S{�����U�]p���b̗�K޷MDq]��F�h/M�}�Ӛ��8)��qj�F�\%I���yn��2��"ذ��Bg���5iŘ���IuP�Q�4��[l��)��(b ko2��Ks6q{�^x����Z�E TcL�"���)��}Q��Uv�fO���Ũܥc=éF� ���[p�����r2�U48����p\�d:�M�"X@j�f�̵�n1���+7�a���Z����W�G=�q^����{5ڒR�^�Fi}�9J���o����o��
� ��SKM{���3*#����d+��*�%W�M]�.�'\���
y/��B+�҆cٙ(-�wlh������6�mN�0R��<p���_q�Ɣ�]8
iH3!ܫ�\�#�b��ցC�O��γ\�a�ѽ��2���T�W5�
�\�����3�ug����Z��L��аbe��R�Q�$QA;~����h�H�cf&��<�{�U�}�]� .��@��7U]�}���F�	f��0��z��i�,��DU= $o���TY��\�+@��7 ��I�o�gI�t���T�� &X����`��D_�7 ���W�X]�NGw�����{$�|�S���E��D��%�O�riB��qV>�M�G���Je�ޣ
�i���G�H?�TW�p��>;]���\��-�o@o��F�f�w_U��bHNǋ�S�s�|� ��Zߝu@�ѱ�4�e��UBNV\����TĔ�
QNY�o2R������ꑾsO��z�+������ߒI�&��1lE��Xw.%�9,�A���@���� �_�G2�}�/�b����������P�4
���L/[�蓷�\)X�sJ!ϴ��~Qk��Oj-�;�q"����F�Uz:j�����H�P�}VV�D���_��rF+d�>��PT�ma᭻B��V�ӈ\���!���^Ƃ�Vd��F���I�������bG1v��ap�ELq���93���s��2R��K��
��T��DٺPp>^���{"��h��};J�'F_'�����#����'���&�;�y�w���R8�f��N�ư�Rۖ�B���:KG�w+�2*�K{�V9k�?ߛ���K:=r�䭇����(i,3���B��T�m��C�T���94~��9�2���_�VĖj-�&����g��ӟY��_���57��lxz>-�QE�[w��q�V��l��-��ju�=���o~Q�)`�z�#�~N\ʤ����VG�~����;i�,�(z�l�L�B=��{}$�v5��8���4E)����/B��;��)��?���\V}3aY#���b�hӦ�9��8��>�I�i�cR�����������ɇyQ�o*���E,a6P ��,>��hV�������l�o�0�*�rBHKQ���+��tE^�)�� ��7a�!ZJ���9= UXa!^Բ���b��h ���JZF�u�3��H@e��'��a �u8C�E|R�%�`D���p��s#
{�!�lY�nE"T�W q?��������dz�NlFͦ��T9�����m�Ϝ�_����:hh�ٚ!+��M
Cf<#a����{����V!'��ε�Z�K�d��ǯBŠ��W���v�,v5c�.�
ۤ1�Z�,��O|��[������]&�ɫqk��O:�/�6�%R�P_��u8�����Amr�'��B��8+���c4�Aۑ��=X)�����w���Ұ�$=ܽ�2~U4)���PL���-I!u�]�8?�~g6� ��(�W�h�E�<�9a��H�f ��])t�҂�@�?�>�ʂ� _�`wb�x>%|�Vɺ�Rw
��U%��m�+<;-�(����l�N��e8�+o`@^L�k�1QE^ҭ��[�C�'�,�y\�#�\���	r�uT�F7�}R�c��8"�t����9���������;��4�}���4��2�(�A����03�p��c瑱З�1a��l��f���bg˶��Q�N��yOH�5���LlEᇟ����*�a�3����x��2���Rc�PV\���&���s3����Hm��8�kG�Y�����6���j�?J tV����ie�ΰ����s���-hlxuz��}aȔCE�G�
�&5�]^��K0O����(�y���غ3�e��5r`���PA��#��p���<\�Iq�mN�*�z�{B�fk�Ƭ�2x�Q`T�f�0�0Pc�_r���ֶ 3���*O��8��/�!Aݩ���"�t5h9u�3=p$e\���nc����u#�x��o����k��G��?����u���ө�-����ceu�ñ��n��E1�XrCK{��x?���<�K�=���fa�ZFu-l��d��^N��S�����ó�ޖ-���2	'�w�`�2�f�gR��3q����ȶH���aw�cQ$�j[L�\��1�mG\��J4o�����3����m$�D|O�Y]��~��|�R�����Ðث�n���+��h��Q3��cp�y� �L��A-�v*�[^�~Ak�&M��ѝl�
��M�&��G��nB��;`�RГ�6�D.���D _�(Mb�u#(�Ȟ:�v)�wb�W���Kd���M�g���4�x��V�~�Q(�+��Q�ܩ�'4�d�=B��*���XEF��Q}ٖ���q��K�tFt��b-�{6�?�m&̀�l<N�X��C�gB�S#p�}�d�"�\6fC�q��U�6�ʺ�Y"�aD#u����64�o�&���\t�f�մ\rt�|�y2>��T-?m�y�S2�{�g"�y̅�c '�S�ྗ�>��}�����X��&�Ta�"}��YB���60��	#N��:Q�o!�?�=T��	������4ULW���j,����t��C��*ti�t�,�˝���{�;�tv�7����C���ΟsT�a�z���1l@�2ԯ����P ^q�1�'ڟ/�⹋* B '
y��Ts�y��J/��@d�O��"��3��
HN�`n������e��,��@���O���J����cX�Y���5Q�������ID��4�Ɇ�`L��6�p�/��B*iE���۱$K9��V�T�MG��q�g5�yY�8�	�QW�,Kr��b|Y�,���Jh&��)�#��$���S(�/T�`�1�E��C���.��[�X�e�Y4f��Lr ��(�Jq<����j���Ղ[#���DE-�l��E=a��î���<4�Kl��H���-���h֑�[�D^� ���o��,�ۓ�vu�a�vI���c�M����p�.���[�|b�)���)���srd��*d���]����W�)G~�|u�W@�_�8݂Q�ǰl��J=5���zf�gB�	�]28q�Azĳx�*�GH��!^ʬ�qf`�LOQY�@Lw���E��	Z�A� ;�W,E<���W�-��P�J`dĀ��=���5���9Uw��F\�!�cq��Q�C�o����7�Tp��k9R;��<�U�ַ_��q�+w�O(�@`ϱ�k�'�4��A���7�e/(�ɾ�m[F��{�_M�~j؎'��c|���5�:�z���=?���[)�r��b1�^b��SoPyÈ��RaՀO�h�߱���u��mD��u	4tf�0�bZ]�o�R��0��� �����V2D�v��u��,���/���H�}E�L�)n�4˼V0>��%�"-`����J�;\��y=��tu������������Y����4{�I��\Td"YGc2��@��n�m�M-#�ԋ�F�aN�Xs��bX��CN��b1�� "<��>y[si�3�h)F'hf�U� �{��Юc�Z-X�9hct R{Jk�8G;����E@U(��G=�i������X,G�*|��(̐y/�cu�8_������|�`����R��(-�V:��?���|�����r��o~#�NJ��׼2&�Q�M�W�\Ϋ.��X��E� �M��MYMk=Q�xvy�JSn"G3L'�H�6o4�N���8�{	�P�;����O̧�#�R���^��ퟄcp4��.�����K�i�bF��#�Q:;��?��8��EN������Kvӻ򧴑[�c���}$��v���-y��*�e��(�iĊbkv��,n,ܓ[\���=����WlX�����%��l�H�l���r�(	�W����yp{n��c'Qp��!॔����
��a1wTA���|���84^m�{�ͯڪ)LK�b��s�C��O,�L*�q&�D)�#T�-�/��`�\0�/2�0�T,�>Z u��o��9�$��'�JN�E�k�VD]�㽙�03a���lW����5S�ϩ"ܰV8�=-<�#��!e����.�|�1��\����8�xA{�};��@[�pI������@��(!�8W$ƌ#�u8*�f�1��Ei��5���`��U[u���.���V ��z�T��|eJje� ���B�k%E+��5��>p�9��僅���_���P}�G���tzZf�3Ql֐(L:��J4(0]�Q�Nnř\��E6R��֙W)�p@���v�[Q��d` �R\���]\��(	NS�G���̘!JU���ܶ��[���n�OE��e9/�T�M9.Jo���Q�j��Ñu%��xT���-?1v�<��� �C�&��u���-���,h(�����
�u��
b�B�K�H7V��±t|m�kg���hL��3i��!@7�|��C_�"�V0�O�Hx�c�\�$ϑm��R�0(5zȔ�r7?�����Җ1R##�'�g��j��@g��k	f+@�Pn��%�~,
��$��#�7oݬ#��A��Q��1 ���iP:�w���IƲ�zћ��$��
�`;���lyĨ�˻�5��Ux���k��v2��@s�-��e|�l�%e��8�Lm���L��vd�ܑt��G~��?�zg��F�Z}ץ��p����VMT%	zT�>Z�EH="�a�Ւ[�s�.�p�:�0/�'~r$ˊ��C��O?�� ����l�%֫m�Y��N�.����������L�	��$�3����7��6>
��@q�Z~b��d�A0�3m(��9�I��i��5�@��^���gW5�����������?I ����C�n$��{Dgķ+���t_|���g ݐ.�˻�����������8Oz���{_��e4w��U7�<~���'#O�����Bu���	ֶR֏�]�A��Kmy	�uDŁí��@R<j:�����۳�{��D�AR;��=�9�h���S5H�=��A�
�{m%��X��R�!�����sdũ������5�j8w�a	�l6���t�u��c7�oqۃ[��P���À��s23�k�_� ���U��	���R�&�h��t?�	�Z�� n�}����
��	%IS*r�PL�W���R���@�joQ>��F�b����Y���o܍v�go�z��M�$��"}�r���ir�֙��3�D�.`WT�w���r�d���l$��5���Z�����l���E�^yM{���*����L��Y]�$EFؕC���EX��h�3�X�ͪ�:a���M�4&(�����W~5����/����Ժ=1�!!�a1Sb�(/��6?_'>�>�$Ўg�Qc�ޤx�*�]m�hN�ֿ��?�N�+��H�[���)JP�V%�b=V�B��Xi���g���!���8�Gԕ�awOj;T��o^J�;��EW�$8�ډ[�Aq;��.RD   ��"��/��9!�|�*}��]���D�!���o2�-�������,8n��r��bG/��: ����.�a�Y!RAFx�y�o"־W��M�y�Q�%657����c��ٵ�����o��Ŗ�|o��� �xP=��ץ4�H&R/��~m|�c^yF��g'�
�vWY�WƎz��hď���jU��^��u����{�},� ���;�N��=�t00�ÁE���j�7�j�|�
�U���,�o+��$��Չ�I~��5���B�u�L+h4ۥ�a�K�P��Dcpk;��~�1��oU]����x�T�Vg��%�
�wh�2���o����|K$B�����O�a+�vW��ƉV� ����	��?F�k�o�h�;`g��@�:[:��Nv������ӓ4��[��
�G(A���`R!� h�秇�K�Y���S�{EH>@�7�%x��1�.4ƹ�2����zj�xȋʡN��e
XB�zn�F�2��iV�T�����H��`�k٭�1��eҍ��2�E5��w9��r�a�(_g"`���S@j�ʽN��p��78�{��CC���?��'8&LBm����^bfV;�H�Ҍ�G+�^ſ8�7XƉ��~��	o���m�y�)N��35rx�]z�@q�t�h�,�%%1&2I.5��o˳U�v2�-|W�h�fS뭓(<��������2hY�h�������0�^1���&:h}�7�Q�eǒn�����5�>|�(�DIby����%�&x;7���<H����b���p��!� z_�Qq\ ڈ9� �����h�%w�}_�*?Ď.A[�ϻ�X8�������e����j��V	�x"����,�P6{��P�t�Vg|�n$�0��I/�@�����>$���f��"N���x1qP+�Lb���u9��u�x��ȃ�M��R9���j��n��Jq{lŁӘV]O2=�bsh3�g�󛱫�-���x,�P2���qW\�	~Z1g�M�2�t���\�/N�\`A�B���b�΅2%�v���3b��hn;�^�R�W'�:���\v�8��:ۛ�,:��v�m�tG�'���0G�W9���%���`J�_�c�o +))xSo"C³[s#߫�o��oɩ�}<c��Am&���gLv����i=�=�����!n��wg�>x4(6H5�4�d���$�U� ,��3�,z�t����}�zC��K���6��@��0B�`�����"���T����£���+�z��ox��C�]�-���0�,G�P�Q�{�+��2��� ��t&�l�ļ�Xޯ�	a���~ƇE�Z��YG}�I^��Mbx�_��y���Cx��h�46����S֒jy8VT�<\�.b�M����:<��Jb&�E0�����/9�xƬ�#���p�N��v�*p�h�≚?�̠��<7T���Z޻R�1�8H�]�Z3K���3��;��wp"|Ԇ'/�@��1t�����e�A�?ں����_)�дd���xf�>3W���\2�3�r$1��e�GN���J�=��S|��[`S�@��s�	������ 5���ưm�*�w���f�Ca���9_	*T��B�qa%�gsҦ��ê6��z-o2�&�o�r�M.܄LݢC٩ v,�Z����L�r�S��lѳeO�Iw�ʲl��Q��z���D�� \@�p�\��R�rD�Z�_��8k�4��<�|I���E�"|����=;Rέ{�ǯ�G�7�ֱ0�.Ƣ����4��wGW�d����i��_���`�o-��?+���jXu��h��ak��� չ	� LT�@i"�a�٬M���_8mk��Z`�7�^n6N�*��ij~��� H�Dn�eT(�x����D�����њ*\B
7]��쾢A�?-�����)�s6��=�0U��ԛ�T�`4u�+�"�"(�[�i�?�a�@_���K�+n��r�/Ҧ%;�ܧY����&c��v�����q����%�j�֜�5L{����6wӛ��$���Gc��S!Q�n�K���s`�J]7d(@U��2�3�+B�a�Erߍ�,\���_�}�O�:�?K�փ#�6�8�\�~�Nm��&��]!.k�w���k��c>�t�Ď��a��/ʧ������W�$T)�Cpj+}]�q?��oP	O�;�[�ew�Sbb���x�'����֤c�y�G*a�ֽ��6��j�*�9~�Z
�m�D�U�a=�ZZ�g� ��:���рsu��!���N�c8ۊ�[�NV$�`����3	'�x��҃]^�
4��(�<Q�͠WBf�X;�]b�w���D��P���k\1h����*�c]r���Z�9���Ş�X�|��u��	qs*��׋c7{����?�v)W�P�S�Tm�x�#��thJ��Rg�N�[oO:��Z,����������o{^:sN�vc�3p	���8�����ۿ�Y�����~T9t&3�ѩL{vd%�!
;�g�?�J�>�9y�#�1SW��~�C�l2'��4'���ѕ���5u��[<MD�qalF��؄�x 5ӂ�� �Xz/ ��ט M�2��K=�4CFD4�^�_yt�,�H�dWS������
ײ,/��4�8������q P(��Y�dc��dp'�ʂc�͉3�f�f��%����s?�����Ø���|��_��G��\����a�[ ��'���ѡ�ӆ���x��%_��R��w�u�%�34>t���d��orL�0lG�>Y8`cێ0��\���DP��őQ��c���1営��-X�1Y���|��;�$���M��W�=+��/�aS%�&�,K��t�֤��r.�=$��c �5�~��i��9i[�&�u�����)���#��
�ڽ�͗,�;Z0�Q{��2NQ���@��05�!�h�ȕ�)
�< �� 0���T��r:p+Ǽ�Z|� C`�rdF�j ��������`nLp
z��j$�}Ƽ�)P8�PI�I���Cn�R� ze��Ev���o��礙��I9��u��g��X`�p��������L�v��@9��cC��s��'h1����9����"����z�����Gٲ�w:����U!xE���Ui$�y�(�0�7�$�3>L�.Ҵ��I&�l"?�9z�T�g>Q����U T6�����h�Ն��\�!�{�)2���%�V<�����l[�f�䢈�H���>�KzOo�,W0x� 9-�1f$� ��vl@���������׃���}���M�����zl�+�Y�Ħ\��S܇(p�����# �)����)� M-k2������_U˸3�a�p�b�#