��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ� �t;l����a�Li�t���A�����������JRs~��Dۍ!J�U�|�4�_OIi���/g�<�˯�_����t}^��[�.�Q�*����,~�R�97��6.��n7Q~%�������)�%����a��˲i9Wԟ!���f��|����W�Qt�H��/u���0��Rd����O�I��y4l��T�B�~��
��ƪ��s�:2����ǆ�������rã�*&���3␾��d�<��n�j�%�wi"��]��[p�m���I'��=A2u5Kb#p+���1�I�o��!K�7u��|�O���2�T6�IL�)h�mE�z�3k)#���G2��:O3�Rk=�r�;6K�0�0���¼uGdޥ_yl�A)��z0��g�b�s�m��*��N)ite�R�P_*� Bf���gQj_���$ޣ4WHF��mN,�Ro�{V���:}{c�h�5�-�$K�T��e��?������݂�����*=
"�o��U���f�M9�J�^�0��?��Ռ�\da�rw}Γ�i��&�Ԓ$�LL�=����iÃY����
ў�/�U<n�c��k���m�Lӷ8���_��x���̐����C���u(��5���%����uǁ��3^Ɏ���A�)�)�j����cP�����E3�����v�62�H�"�e���bA�G�z�MD��}�f[?����iE=��W���l��䖿y�c\�D�
���%��([��-��z*6FԮwƱ/V�Ơ9F�d}I��S����#g�ιU��r�VT�!�α�N���7gU�-���K�lm����c��oi!v�!{����٫r���_��@8�e��+��V�Va��6�~hK⹷k����ED� D#�L<��O�1'�+p]��]T�̋�NC��Mqh����(X���u!h�m����c�)�w?Wt�	Xe�f������Z���i7�q)#*�=���o�6�pݸ��� t�1>+>�Bl/��|̵�+�gw��b��3k�N�T,�L.�f��@��A�:�Th�,0S�Y�Q'�R�� ��0~lr5�Q4��� >b�T7���}��,�O�Ǎ��!/�w"N����6��]S���%�*A�������T�*D�5g�p��rh���\(�4���������ϴ�*N���f��J3� ��	~�dd9VN:�#�5t��hM{YP$���#�f��ESv�tJ�χ�li|u(�
9�`��請�|�iئ6p;�J��l�xo��U�#�E��_���"�Ց��Q�IHu�L�|��Ut*GiQ��m ��H����:��TA7?B'��](7xa���T`�/���/kJy�>��/k�'�Sx[��F���!'�k^[P!�����Eo�צ�44W�4:�GD\�+�<v̰�c��YT�2��D�����|g��	�.�;Ee9: ��3�V	v��ӝp{���0")�)�<B�N.j�DT�Q*��Ծ�1p���luB�,h��Zh�]��D��j���a�o�3bZhB�G� C���
�H�M#���a��[�C�do�(�$ �;H	��Y9Ux�J�YM,`��O�j������J�A�w�c<���x�h�Kt􂛫p��Eb��~d�ZۯoR\���;��yhsR7Z��'=�Ǫߖl����Cӯ�����d��m}��#C#��N���S�@�?����	���9���U3z	b�-��i����5����k��4�"x���w2`�^غ>������]=��$D��k!����\ϵuzy�z�' �hx
��JP�c\�b߬��t4E��?�����Fz<�"�<�pd�y)��L�O���'Mu��^4޺�V����)k���%S�:Fw_���0�r@6�ټ����φ� ����q��X�N���	�1-��y� �p����6Ɩ^��| ���m��5���Q���K�Pw7�0'�����tz'6�>���;Z��m����M�wk5�`c��WzF��W�!�X�΁\��0}���7O����|��&���
��'�Hi�Di��U�q,�"]�8��@"41M��!������	ɡ	��ٶ���HJ��Q��ʅPnn��=bd�}���Ƶ�q�.���R��W����*_:+�a�����~qǤ��bQ�M2�B�a�>�k>ߘ�86��Vƅӥ��hU��@�W�N�h�[G����g>���N"�ӆ����t�⧰+w��  R���,�3�C��{�w���tC����WM$��./x
=�>�~��.�7~B��#��6��u�4����a;> �B���ϵO����Ng��Y��6�^��4�:���F�CC] .}�1�j��L�H�Hy��$=�۫l��s�t!�;��Y�bIo��,��d���^�J�����A���gⲿ^��N����6'�oZ1HXC�X̸�G� �}�"}K ?�\4��M�(��G�s�2�h��F��{"_m�;��М <t��r=�d�����ʺ8%�'�f1&*�<{$��	E�hb�^���%���NoH�c+�dE�U�*���� ��h+)�,�� �ib�Fí���QX]��v�j�4�UG�}�M����_�k�v���5����,�0�.���=
�0G�a�\��FE|ʈ�D���d+7! ��h7��:��,��kݭ�ۭSc��å�w�4�IK��k�;7T�A�j�v�d8v��3�sZ(�'
���@��¶�cl�����d���1t>Q[ƃ�~6���iD�̣�rM,[�7� ��8n˪,&�5!����]�}��R���4�qw��*�C`�s��p��I���F����6�d}��2���z�%���3��*5ո�k�4/G�$Kr-K2�Qڋ*�2� ��T�1��Ab28�z�up���D �[I��R��׹X��� Օ�Ė�~�&. Zz�U�a��K�k��!�A
Gq���䪹"=^��j�x�0ɬr�Qq�yv�@�w��F�&�'>F�_���jN�ʵ]�4�,p����������K��u�D����| B��&���a���c4��fs^���Kn���u=}�`��ae�=�L'E�H<��A������4�E
��b�`c�&��_��'N%�_Q���<��Ns�g�rr�Ua��A���?� G���]�]���P�>h1���c[�@:��!H�4��zl�s�+�*+>{��i���EV?�*����w�'�`@�C|��/�o��#���.91�)׸���6_�r��x�0Xc�6���*��hIJ� "�,\����rk*@LP����|��$�>�
�����U�Z�ˈ$�@�bi'��%Jx&�wG4Yąי��uՑ+�bW���bx|����32�%2�L���6s��\�X�DmXr$)M�:n��z�&�}�Ɨ�7���uG�{��KC����e��Ӫw�ef��~�n�"���r9~1<0?�7?$0���[��;�\(QL��<�"�M�6����aL�A}�����\�+���,��	"�1	���G���'����$����^l��"0�=�0+z�۞}�^Âp���ۧ�8�O2���k�����Q����������B?���%�̲��Y!��;����ZF�o;� 4�vAb�2�JI3TAn�,MI��Z�[���:�^��L,�a��N��M+����is��ok[ok���`�:�]�[:-<��c�o7.�cV#4;Eպ���z
N����vT��欠��I�p��0)Q�H|�G���6��Lbɴ�?	 N-���8�����߮��Uzƈ����58�	���D����s2�5���Xh�M�#VQ�xo"f�l�q5�=��rG�c�"��[��Ԣ������ܜQ����,+0Kv{@E�ҦX�}k�َ����IB��F�����ѺډmՌ��iC��*� �_# V��f�Hd�����`Xx�k�΂��I+
�F8�?���>�6��-�L���owi����]|����@՘~ɉ�)6��
����9>�;��wG�ŋ=D�}1Ϳ��:HB�/rG�o��_D�j����#�~�f��Ŵ'Ħ�9(-�o�Ĉ�&�T��ai��T6ɞ�#���S�;��7,:S �r,�8��㜠8������{E�/�ݾҒ�v\/��͟�p����������g|��=�۬;�o	z��<����ic�ǻ�>/@/q}�[f������8�vbz�G�mr��#Iy���w؟�=��ο���4�9��En����fQ�z%@��	XS��v8��=�Lꙣ@� �`V|�G���������u	O'�����g�y1��ּ��ok]O���xk����ȏo�X����ߏ����9#J��p���%,�@p�Ĕ��.��h��jɦxx�� 5�쵆��?�سo�~�D��RCҿ�3�~�׉H�JF8���;dj�g�Q����`̉Yd�\�E{
,�Yc��uLLa���e�!K05��k�^P3��j�"�Dލ{��]�`9�M�`>R�b���9C�������9���_v�FX�'�&m�'yS�]��nB"���Я������I����
�S�(ge��i���Xj�R;O?1�S��h'���H���a����"N�K3R��41suw��J����,ǫy���A�8�l��all�`�j>!bs�	3C7��è��ӣ�����x�n�r w�H�A����u��QX
��%�E]��JS �}��K�'��3�̊�߰��p����`�S��l����/���4����^�@ѭ��,��W	�Gt)��3��n]�u^Ku�:��W�D��L�,y���Q��GpǾx�(X�P�'Sx�E��&u�O�D����=��l
̇i)��1g�ʭ��g=���R&�����R�s6̭���(�[�p)�`d�d�
-8�I����`e&2�Z�?_)�_W�#�T挐W�}���:L�6;Ìu�T���-b�����;�OA=��g���x��{H�!�$�S綊��Ф�n�n!����RL�� &%�Y�D}!'t�q�D�}�dv�CKp�^��dκ�����F��{�����^���v��I�|[CE��n��h`J�+�>��Hn�n(C v�Oʨ�~��~r$Y �<i�����j���zU,C�w��3��Ɉ�'p.�HSUe��!�$������)��5,k����Ш'�����oa��Q���"� ��G�����`,���R�D��p�
-�j�@��u?"����v+�9e�\�b�;��G��|�P2���{��RW:�
�TJ�.��A�z��* u�Z�=��;ڣB����B��h`�(5N�1n���
���0.aߑeoU=�í7Bd`bk?���n�0����9�H6���Rw0�6�ݿ�;�L��sPC�KB���M0m�G)���5��gr�������j�'^��T7�ψu/��+-�&x�2=��aZ�%���=4\�O`�u�,���޴��8���?ί6G$���b�-P�s*�`�j�����|���
|d!��gΚ�[�Ux�93�b��:��"Lnğ7kb�鷲7 5ߩ�?���m�7��|PY*e�����D�y��kLEq�s�n^�)��/��a�k���b:(g9V��+s�ֈ�)rl��0��m&�n��Y�#:=�WV����C��f��3��ߨ��y|���{WV��`�b�r�H��R��n/�3��{_B�oT�A��6S�2ca=w���ŵ��صz"Q� ��'tl{&�*ƥ�D�F?oON� B���R*�l��;�ќ��䐸��"K;q7�!��&W�1W���q�u��p�0!0����y��v�.�*���2���A>���Lr'�x�qLS=�l��:��_?�z�ThO��`��|�Ʊɜ0D�Ë��	Q߫�d������J����F�$0i�Eqi��$�aD��m:�m�r�sQGs��^��TX�r�.���*���3'��g��5Ag_[\ Q�,`�U��,�m�?�D[��4��0�����\��4�n����f��l*��0�Q�~����ȯ��J��j�Y�L*��V�9���!�
�J�ٳ}fa�YL�p�E</��>K��(�e���ZV��ĵx�CQ�5��[�܏�?ʟ!�_R�m�����"��� �3~Ժ��1�:ܡ��E.h.oa�A>�L"�g#. ��t鎧U��<�T5�}�y
{Z[]M�Z@��zi\G�~������t�e2���Ω����bF��O�wh�vB��]�*�Ḭ��	�Ww�z��t�J�.�����r�ļ�u;>sG�AK�/�7�37�>�0=��^�����	Ҋ��Ҷ�����5�m���l	IW��{��!��������Z�F�zP���3�U��g��1Nᰃkd D�5�J�X�?��7'��~�~�-ܫ�c�&��s,�G��g8��@�;��m9�@�r:�,���*�54��f X�l���K�S%S���E	<;!�dUce���2�\]mm�����-��NuD���-��IҢ.Z����4��}�E�����)���έI6#,	z3��~�ס��WL������K�w�2��{�t�Ae�j�r1DB$Ϗb����I:D1;mR��ɣ>��%�������gj��a�O��m�ߌO��{���~)�0pe����P�qɃϹ���b��G�O�(��rhV�vcv�DV_����	��݌1 eŲ$��"N�DkG5���ЏWB�O���?k
�O}�t�k@��U�G �(9��#Ы>txl!em8g�ߗ�J��D9�`kH�U��}l�R"^mj.Q3����4D�ɘ��� <S������58�aHҲ�Z�J%��a��C��AD�}���2@=��s?'�y�5�e����B"!En�yS+�����bk�2G�e�ŷ	��2��XEGπ��"�|)J�P��lyY�6<��O��o���1�p����c��P�a���R�O%�\�6�P	���Z�XA�f{g�����ؐ��]�qs�4��`�j�Ñ�>K��1&�j�:U�jR	{͛�
������}��*l�*YlÙ� 	Ņ�ŧ�����2I����iN̐or�~Q�4�)��1v�=�����R&'���ž�aKJ4�젱q�i���b�wL5��`��w��3���%N���'��_�Mr����{t��wc,E=1�3n�<�4�Rʣ�L�yG���4��O�(g|�Ux� l��?�?�3���������.��!¼1q����1�����o�;"4�0��`��.6mt^�%��ʣ�T^��m`+�$P�R^�%�7�H֥��6nʊx.�uOp�SFK���(ݱ��+��\��*�O��D��ϋ-%虽�k�q�ұ�	'���	�`|���s�������S&���8��Vs�)�T8�]>B�b�j�v��?�R1=Ds`0+:������b�rD`)�g��%+a��2G;f�������^��K����	!jq�m��i�u�cw���q��]o�0�6�)�v2� �FA����s�V���Ғ(K+<�arLS�*���a����~��,�˞��Z_q�p_��A�P�r��TFv5M�x"�c�ő؝G�I��5���r�M�3޿���������I�M���0��֖�:�e�R�}I�����e
|D�X��7�_ �L���+�V��4�����|#��ym@D��)�'��Po���o��6"�a���RT�|��[1�sT���e%e-ͱ�[Ip��%�IOjX�N	�B2����^JZ�Ț�����y?u&V�T��F�?�l�y�6|r�K���ē���E��z���}��֦r��"p��|"�qմ������~�*�pOz���j��4n�^�S���
�VЕ���۶3�j_�s�G�n�b���xˢ}9�/�����gf6N[S��w[p��g��aC�����(�PMQ
չQ�[�~�~ d*.fɅLT9�`/�<#�����o�Ԙ!���Z��*��]Ǔ�5�=0y@�o�������2�E�UH�j��_ި\q�ԿH�!�z���6=�
nc1"T�9ɹ�����8iUh�:F�<��t�'@�S8\(.�/tF�}|�g�� �<�N4�ө���ґ��r8t�?zǥh �,�>��ܘi �Q�^���g�ŴQ�®^�Z�T�m?<���߾�h�E\���	R�B���?�����p�'�8�G��)ڃ���Is�NG7��D��1��$�a��FU�4c�m�jt�R��6��xV��%ټX�� Ī�{�D[�K'���	�E<Wdɒ"u�F�{���s��B�/��Y� �.*���o�o���@n&����X<�o����)�GXI�����(*��0�f.�8�+��|i���o�ވ�E^���h�41�}���au�ʟO����Bt�LK@%��q��X#�jH%����y��y���$EO��H�<�Щ�n>?2����(t�|vqb��h9��0��p�$z��e��v��;����L���U����P0é%]�fA��đ4��X�{*)�B/�xJԹ��Nn��{��Z�>}��_��}��uk����{-hjLH��L�1��f�Z�>\N�����0�L ;�gQ�a�
>C�(���smr�A��P��7�u���b�W�Τ|�� �q0N����պ��|�_m�I���J�g�u�*|�^���S�F[b=&7]�^�E����^�$�������xX�Eb�:��C?X4���q���h�垺~����������U*͂~|�!.���MSL�0]x��.�J��P�i?�MZ�M�*b˅�7̸Y�,q,����' ��1��v
l�%K�Lhd�N��m�Ǯ?ឬyc�x�7 ᭮L�q��4��̎գt�9� k��F5Ql�N4 `b�J��}���XŌdrF���i����-:�L�ž[,�O��o� n��Ҍ��"	��J�A�:�t~a7v�!��,W[Ю69^>�u+&'F�9�����o�Ǉ��@u�HK+Ǹ�[*��̗�%����;����/m����⩊�P�/buٿ�%��<��""F�d�q�ԉ��r9������9��S�g.�w ��S����[�waj�#�o�鍋յRK�E�U
���ҥ��o�jf� b���Xs���e��,y#�]����F��/Tᢤ�d���ݒnSH)�
�jF�"Ն%!'V�5��`oU��`���r�!?�Մ4� �H�8kr�yo��!a��LIvk�7����~-8z�Ѡ�\�U#Π���U�@)/P�U���$�[�+(Y:�s ���~��*���u��{�R��4i?%���뛔��"V��!^}�O͸[=u��t�6�B-�HY��o�f�Oɴc��p���G�s�,����y���|��|��텫�^�U	�ʙ��<����h��?��|�};Ӽ�#�L�|��XH���H����ԁ�2�������b��$/�*��\��N�~��q/\�d�	����W�Z�6��o�*9�ڊ$>i'	
�*��gf+���Jފ� ]#�@�@%S�y�뇎˹-�7��*���<��#|]>(S�F��9a��O18�";��NY�y��h0_��������qo�lHZ {��i�~��
�X����Z�O㗢��c�H�6W���b'����[[kP�~��Ӂ7S-+Ļ�L�U�r'��A��swa���p�/Ms�Ϩ����&i}�o�+L ��/�C!�/|S�����w��40��o��7�
}����$���E��|�������2�%�����겑C��F�Y�I
G���W�􊶥V�ȘJGM�W��(�'B~������\9|��ZX�%S�~���]��|9!��v�h���G�A�ٸ\}?�ץc�5D�W���z�}F&�/� +������R�������mY4(!q<qD�-�1Y�쟤�q���'[�ĜD�GS��� +6(7��Q�:�oy�1���x�5�)�
�`�Ge���s��:ꦠF5�,��PsGj����\��Dӡ]��h�f?�t/*���i��ϖ��Sv��/���)����B�p�T���	f�FutU�j����t:��Z��(G�x���3��ܥ�+����v]*��g��^o*x�G�@�~i�j-�BBvMڥ`��w"�
�]$~�^��_����f�)�R��POH���J�u�`ȷ-�����A���1�^
$��}��:��H�Yӳ�w����)�*���<���e�Vd�G��lz�k���EL' %
y�x�^�%y=,���X(�L�&3R��F���z��+�V���݇Q�ET�',e&
�<��ی���Ax:L��$x����/����J������D�?�M�gP%��^$�F�#�P(�M��� ��%m���4���é	S���u`�8/<ϭ�� �7P����)t���o	,V�FP�k]C���`���t8��;��=��y*�\Im��AF�$����7�q�<osI�*�����(R�$>��f���G�R����[�o�#���C�v��7��lJ��`�Q��i��hה��݉%�)�Y]Z���[U$�BI>�~�+48���S`��+��"��-�����)�����D*�:�Ц���U<}MhG<]ſJ���%����suٙs^��{��3^lO�@x\x�jBaB���E0I��н��|gu�6[�EŪ,7�N�j}��h}@�Au�6(x�q�#�t�~A w��]]tã�hR�[�i�\�oQ�,9�[��0�m��3Y���m���FH��%Nb>*���D�e����0S��-'�1����ӽ4��K5�+m��oI+�[K����S3J{��?a������%�>�[ù%I�k\3�e���U��#>e؈�M\����i�P����Z2��k�}��a.� ����O�2�A(!�Q��?���<������♿b�6ߚX=�����@�B#�.g�CF@%{�7�����U�M`*��G�:R.�Ӎ�՚���3C�[f�`R�"���~)P��/c�G��P�3�nZ��>@`v2����92�*���A�@4�R&��+�]`jq_��X%�����f�:<K��JށιVlP�B��x��fDZ��Nڊ�6��2�Z�L�Ť�Ӧ��;� 鍺���?@&A/��ʄC�W�[Pe��6f��?%��S �Tm���6���X���Z��J�ټ�NNdr�z�	����S�y>7J���0��y%��و
�pK���P3�� i��]U,���f���Z��$�GR)���*��[��4��^ʨ��Tl-� {���{!�ؘ-b c�T%�X�A��6h��G�Z?1�`u2 �S�qIlh���	*��c��S��Y�Ŧ1@j�/�h��|��Rj�_^�/��:3umk�#��j���}�)�3xm97f���[�W3>~�2a�{o��<�E~�m�MP��/�_e�A�S��<-�#����Ko�N����B�P�՛)a�
'�;�Ðu.p���A���9	�G�vI�+�R)G@����sF�j��/*GujI����#�H�ܚ��e'�	��:,9����|�c��d7`(WgFW�Q���B
�:/��b�X�Dj�yN���B�SbJY:��J�l+`eA����U��0ʫ�,|9�b�l�X6M���~ሸ��kĂ47"Ÿc��=�_b�s��h����'>��1^���='��Y�f��[�(<���N^k,Җ�K]���@���\�l��>��؊<#�o��
�J�q��R����&�ga��z�&�����.�[֐C?�W�l�"N�����:^)�� 1r�����QG�W����iQ���rb�|[b�e�槐��2��/^(�$ó�:z5e4n���Ͼ�(�8S��ʗ2��Vl�,.E%�ڶt=Ɲ�3-s�c�,�,Y�C-��_�n�@�J�g�]@ ��]B�,�S,;<o���[�dŰ�Ծ?��-�}䬦T��l�~EP�ܓZ��~}k��V(�b����Ji�(Q�	�{4���e')2蒝�Mؗ���L�����f<�ib�/��Te00s��\~79�+�H�Ʈ}���P��#CpCv���.�����ŏù7�jٽ�D���
��7��r�Qu�� �l��R�%��Ɖb2�M�8) ����b#)����M������-��rƺ��Ao`���#�~	ɟ��z�;+�!kj�&��û�*���Q���/���s�O�q�V�I��y����[S���/��<͏_q,�J��t<K·��4�dd+��s�u���Y����u��GH�=_RżI7@�^�/Sy��Ⱦ���c�.��e�,��a�(�! 	O ��}?\pfAu�+p���MN~�ɠ�/��4ux�TS���.ln�)������/�B�b=�Έ����&憒Ŝײ�m
z�g�-�Vt������~�5�c��WNdወ�0�!+#_{8�B3)����
�];L�e�k���x"���*��?�G�g/�;�����֙�i�}����ZpB�����U>g���M9<�=��XW�U�X�ͤ�H`(-R�8���	@.ٟh���$� 7傳�+�Z�L���7���Lh���X�&QA#�����Q�fb5����S��XB��)Ř�g�-�,�o�h�O���յID!�E��#yڦxY��)�I��CYXw��,���"�ʊBz��?�?d�D��h��QA�)+^�?��1�����5zbyQ!��Wy��
�'i;��xb�!=���
��$�����J�$��X �AI.�{�;"��#!�F�����#����^��у"��S��l�)���2��*�a">T�F���w������`��/�Y�\4�^ʮ�F(�sX?�C�{LA+.�dc�Ǵ*��A���h�"	��R���o���aI,�'
jt���x�,�@'R~���N�.�dg��+#B�q�
DL�T�oa�64��A�N�d'�q�nN΀d�]��%����Qᕑ����q����o!/+�����;��E%VF�ߣR�"xe!�_���A�J��U�L�6�zW��m���A�k�����t�ϼ|W�Չ2O�#]��neT�My��-��=8����u:uI�:���$�*�y�� Җ��'���0 �y��ķa%���wK��!�)�gu_q����7���O>�zl��fgSf���ٚ�U&�/P��[�ȼjV����a��c��Ԥ�YTqep_��������/�˪;���QUM���^b"/��5\��&rkC�뺸Iڿ��dh,+�߹j��o����H��/
"����y�����C�9�1`���)�kH%PZ�%��ِ۠eD\%��ex ��wvC����^ʋ&BF���*�)���nHP�X�AµqN��X�����x
�����k/>3��wz�c�ij7����I�?x؁#�nV�ϋArɩ�+_U�O&��҈��A\�DD�p�.��� ���៰������H��J�s#�q�.��Rm�Q.}����]g�������|�5������>��M[��o�{g�05�+9�sv;O�r����=�F=]���/���}D��>����;`�w���Bf}T�JQ��Z�f�q�Zt��4E�m;�v�q"�z )�9� Ax�G��p|�:Q1�)K�������yi��lq�8ya/'�����z��a"�>��}�_��d�x�d�E!���ƴ��L�Sp�^'��#�,OMd:�v�7�u�.y$ؔUޘG�3����T���z��ܘI�pe���}^���#P
�Q1�-/�.�`�n�v�@@\x)�jݿ24O��Α�IVu���?4��.F،�4��?r�{�[B���fO�-���>[I�Y��6ɳ��q�=i&�G���DHrSfr��G�ԅ�Yx����pyE��7��L~�Ռ�惻
+�F�I�1����9�Q6�k/��N�E�*���[]pqdgNd5f�*�)/@���`�9��0��7��r�3�%�)\�DB��*9^��EU}g�0l!�>����Г���Vܧ��_zjNP���н~��6�����(o����)�v���?}�5�W
�Weբ`���I�>���Ղ�9���6�\n���.dؐ趒��������$*��meS+����au�bY�p��oJd���5U
ݦ��.�z�ȫRe8���-�j4^�{3�7�crG����3�>�sn���DwV_�#e�c%;�� Ŷ������O;_���%��?��1Bz��M�Hk�X�Ę1��"j!M���ݤ,�z���;�{en~B�O����	�Vd�ō�6���d\���)PUN�Y�F��=�ʱ�̋���k_�`��O{[�7�)�,�]r���pp�fF�S~wm�D��5ܗ�͔�A(�/�'5��qQ���;�%5���|M�\�~��D�[����ꪮ���7�F����&�J[$�-�|�m�7ɳj����sO�#(��V�Qm.���Iȇѝz�H�Z3�>O�ѓ�N���o�Y��[���b@�.}(6�!Z+�s���������UP��:����9��:�E1N���r�R�C옒���^*At<G�2���^�=Hr�I����ҜO�x����"�`Q��ĠDPɻ|��� �h����MSy�m�� ���M6��Tؖ+E_�e˲����e�Һ��,�잚Z�����z�܄%z!�u��O7���� q��󭃠t�p=��A(�9������B���)��H����� q�0�D���&;�o������<B���p��c�!�H�ۻ����iK��XLw��+c]a�1ɴm��C�g�I��l1a�U�IU���Hkd�	��i�x�� 8xJ�*��g����J�vfo@]��(��I�}}Ɲ���(��&���K�y�?��F����':���5O60eд��(�*�p���$�6�����@�K���~���sbcc�s��vɲ#s6���yM���������!�B03jo��P�f�!wx;�/�;���.�j�>>.��a�8&�e
>N�Aj鈭
���`}����6~��?���1�N���D�c�)�}���������!�wu���>>�Ir�ɯU�|�#�E�a�(�{�n����N(�/H'gXk��ȷa
�1l ڽqZ��V�ћ v �e�	k'�/P�t��wvn�8g��'sZ��N{W��Y���������u!(�'i�]��Y��DA��Ì J}�n$����L���|䅤#����L&2�	�:Ɋ���'��?È�\�HI{��mN��ע3�y*D#5��R`�pݮ8���r��M�@�%ˢ����]Ԃ��K��4����>y��[��3*�ph����7!�."_9����H@3����w��Gd�`~��^�M�,@qG���s�RgnT�zt�?}o�X�Q������8�'�o���w��[����z��wg>��)��'�iB(>���ս�$���?���R�[$�����0�袶
�2��=�����{���PTOv ����ڻ6�>��@/k��&�V�W���`�"�/A ��D0���ϺI��~���xq�o��RA<��� ��nNF��C
��/�ڋЀT�9����3e*j���D�]2�� ��)�����<~�P�`l��#�l�y���4���|�VO7��T�0�OO׌=�|m�A��Gϝܼ���/R�-���L�v��ۂ��o��c0>�A�D�)��ԁx�_ۭ�W)-v6�41��)���)�ʣ��av+�V�j�򣁱��ؗ�f48B�˞�$8!�}l���@$w��q�r��	��iZ"4�'��Tڰeն*�,��Ѳ�����|~��P|-^'
K`%L�xU����5j��(>QO	�؉+�2�"�2�4�~N��ʫL�d��E^KWB�[�d������#��ʀ�[�mih�I�q�ʅ�V����?t@qf�DWyY��3����+e�搽�O����F���q� G���Y���U7j��KyK�Ο���}gr��bj�W���8	y��ec�� ��#A//��A��5*�;�I�YJ�7���w�=�h}�|��"oK&����l�7j���>Z	c�w�H&��0�aB� |w�z�������=��!l䲰佈�m��'��9Ƕ�g�2DF���u%k�|�C��7O$�Ih4[�ǣ�\���ָ������y$�m��w�W�Y)\H�#hdipM��g+q�wFR����uM�b<X�0b���~
;}�i�R̐�/0��(U����T��Tb�W��R:3xK�+��E�0�u��F��n�h�T���;�f+�@�Dp<P�%�Nt�#獱u�ȃ���by�`�4��ğ�H+���=_ ���Qb� ��!iV�,����ITþ�vƁ9VCl�0����%���C>��y�%LZ>bA4�q��x�I�
'C�9�� 0��@�!�ts3&� 1��by���$������D3|���f��ڝ���8'C�F58?ў��<�}�2$����"�?���V�b��N �Y���~v���O�V�N���gw���%S��ie�� �����f����Y������S�A���li�HHK��(���[
�ǡ����Z>F h���%�m7���:c�3�\=,L�$BN�8�����Q��@�������h���F=��s�X��Q���^�=ٱ�~����<������t�v���~��K����Q?F�D9�m�X�k����v���ù �&�a+D����i�� ��*Bݻ���S$>p_�����W2�y��p�LX!!z��Rp��M$��1�D�=�D�׼m#��$�*���s9-����P+�M�0����jǃ�����4���Յ�^���Ek��]Z(]�O���=��.ߞl���"x]�e�p������ǻYf@��*��$��5��^LlǄ��i}9Q%�����Z<�Z/�v^P[M����*�>hwZ�Pdy�1:��x�����9`����ʶ6�G�[�M0�9s3�����	���~�a�9��|>KV�^��m+���WT] �z��$�7!��xL��D �1��@�ػ+;R�'vfT1��$���e9#6G�c���g�''�;�����}�#*H���b�Vq.���Xa���a\A$�C!�qz��s��Q�D��O��p�K*��pT�oa5���ŔQ�l�L�Sg�0DH*�F�&J����Â������_P�>+#���\ʐ��eޡ�:����J<����}sW��\��2��T����28-+!̖@ �*ӧ��H�뭱�(�<�d_%n��Q"�ڤ��2�ZEu怏�e�6��:�ԅ���G��)yM��?�:����;ju����+#�-*@QT�U��7k��0�����(��wl��b7���kez/e\l���; 6�;|����<�g��Mߔ��Qu�`���<�I����2���ۡ��<��¼�4����.�;1��{�1J�:F���Y�4g�q�\���r��-�R�y���JI����5{t\h��h)��b�(����,'T����݊?��v���1�D�k�yJ\�X������l��M�W��3lN6\��0��N�N������Lw@q����,Z�2�Y~m�O�=k�^�{�w�Y�KS�ဆ7 FF����!+&?��>���p�\�\�׮y���B�cd�jn�b�3�6CO�0\K��p*���XL�T}WT��=b��m'��m]G�hv��VR� Z|җ�L���Wn�24�1~O����&��}�3+L��#˗��iq�Z�@`��z?�@��K(&�L��Z�"�'��f�򌾱9��*�VO=���À���D ��"4�ȯ�^
d�]���RO��g��!@A��K��c��N����*7�Ʊ�[�'�~��B�V����(��/Np����Č[�Ȟ"�ױ��wɅ<~1�b7pe
'�qm�e|YP�#���Vʿ.U�MEۡ�M"�7ס��x����Ã�Y�$���S�rګAߋ�ݲ8M��cz���o4��P������_.,¢��2w��vC��
�&;=iu(v����J��sZB�b��K�8~Ǹ<�9Id�N�o�8c �<�uGK���vTC/{O�Ec��j*��]��%6A^��sn�1g��P��1�A��>;\0�Wp}c��S >����Xn��j`L)����uӺ<�迢`�X{=��.�oI�5�!�0.�3�ĝ��V��W\5��qgϞ����$h��S���#��n�҃m���]ƿ9o�4�����o�3[@���T����f=�Ta�Ŭ{q���d�w	�e������%�4��P�����s!s"׷e� a��Da<Z��r<sC�k��0/ٟ����j(K���A���5l�& �#��tcM����r�R[�M$�YEC֖�n�A���7�M�����0C���p�Z��X�ٵo�#��h��0��nH e���b9����,��R~�	���XJ�ec�+{��jy��\:@HZ�]�HZX�v�'U�t*"[���j��|1���l�ٷ��� ���M{B6,B�,���2B̿K�F��e���dxģ�V�̂i�[G_e	��M�����⻹����q3�#��3q����0
�7v��mg<�9��jǞ��y��;:�#�@wP����qr7��YÙ�Jێ�.��@�hi����j�U��p��X�����	>��ج���)No�_:���\�����D��Nh�02Ԋ�Wi��$��m).p(o���
X.8��O�6u�2�����Nf0pq�1��|�������%����s��@���~�#8@����g�!�爊�\�H���-��S/����疣4��d���ڿ������T9�yM��u�F#���ѰSiY0vս���+���gœ('$J#~��)ĸ��3f������e���Z��,���/�šD�d��%��1��޼5P�;���bM��kQ$j��✇&�P�����2��_t0k���2�k!�� �_h�h$����y9�Z���mCͪ �	r�h�8Y������i@���j2�v�!�1��� 4������ǝho*�4OҮ@��yL<I��X����&Z�_Ib��ɣ�y��	&�flHY#�Ě�Qؓ�3�a���[n��3=�����}�ܬi��x�^/�������G�X�d�k�&)%�:�:n���is�"��}a8ʖ�x7f��������o*Ex����D����|�sX]��{�.���KA
�&�@��IbVB�|q���o�#���C[��7u;C�c7j��My����v�3��"b�9�SM�)`�=��&���=H���Н���L���0�_Vm�s֚�	6i�uf�g���A���gWR#���GP����%���|�7I%'�['�ý�����M���F�ωe�7�<�B&��\Z`
W�Jκ���17��XRL�}5�"uu�(l��������v���
��8wV8F��~�T0oꖆ@&f�/�x�f�j��q^%���"5΢@�V�f�6�W����cMj��9�~�O;`���Lh��H���cJ2s}�:>�)m�/F�7}��Q4E���F=��\Gk��m�}��0���u���dP.�9`<w?!L)ϳ~F|D���7_A�f(P����vH��n����M�Uj�b�,��z��7����87f�|���_���z�3~�x�1�$`ɣ��q��R%`�\����e~{�";�KPX
Ukd��0Vy��#���#��c�ܝ0�;����8�����y�����|�G`3��U�׶�f�cxDm�`�?� ��Y[ۺ5]�3Q�;@����BRL6�E���7���=��lM8��K*�.@kV��ğN=X���<'���+8���Qh�g�����P�7&�U����ob<a�E�w�=�rV�,��4ck,3,��l�sa��p*�/� h�;Q(�k���x$�#c�7��` ���P�㨎иI�Œ*\���[~=d�x���-�$���9)-\�븂y��F�dG�5�ȍ��=Z����؁���qH謩}�e�G�T�v����60�!	�8yJ����ޙS(߹;�P��&U����k�_1�*QX�XY�&��?m�Y�T~V��sTJ�:�
'��E(�ڶ̇sgY]�Z� 2~����u+��0��{]D�|��Ϩ��}�����'y2����%��6qc�Z�4������?mqn��1�^vq����^n ;����bG�S�۪�X�?K\��t�!WA[>�QQ*R�],�� *CN��陳9��*9o�:
��"��4�J�4�'<@-��Q^���S���i~@�mt�����	�&/T\��a�Y���n!\���C�v8��^2�Ɖ����Q�:b�QfOҰ���T?��J5ه���tP4���?C��<x�;$��-gA2"ͯ?���qp�u��/D�Z)�}D���Y��ܑ˹��=1"�4xG���x\���tR?�0�1�v"�6�����L�������_.�`���}xث#�ʛ�tZ&�Q�R�FsƟ'��a�k�y��Ƈ�`h����D豄I G�J&p�����{ vr+ᣩ�	�0������C$'Hl[��"߱�@^�dݤH�%a��u��b��F�	� ?-_s�1�:/�9�1c�ml6`�S�����	��uW��rM���`��\Q���Rzc������R�U��9K�~[�qVt��:���iF��6�C?	�[˰��A��a�5=�'S���`��|�R�ۅ��a຅����wX���}���B-��%c�ӟ�x3w"�������~����.Q�{�^;θ:���;G�lp���I���5l}b&�	]p��Q���O�:0�'*+�:p�.uOրҒq��Q-��ߓ����+X�t��Af��rAl���Oݽ���ݔ���d��`'��������I��t[G�Qtr��K%�{Yq�9_ �~G%�X�e,bE����#fđ�y Kt�Nr�Og`�nhaP���#��;����d�w�&�.WU;&'�Ya�l�R,����9Ś5�چ���pX�j�~e8��p@j��������k�	ki�Gͷ�Le�
���p�k� ���ۄŎ��n�a��g��s��FК$� ��^;���e��i��uT��%2���h�d(H��v$W.a8�W!	@�M��4��X�h�^�/�M�:�;5��n�6��}P�_$����M��;x��0w�L��z1�d� T���o��9>�����l+L��T�0қ��k�<.?-a���[ђ�!U�NKPd��Ϝ+w�������	�]�mw��V$E��9OM��h��,e�H�ņ��M�9�:E�'KAb��)�L�Ք�}W��EC?V���p���r�f��X����ۍcxm�z[��%���P�.�G��@0tuӯo���=о��T�b�=��@�4�ۛ�	o~�`~��4Jڶ�q�޳���#� ��+�$3��\ ZbTݹ�&^����V%&���xF�c���7�u���&s|)s�787@���W�͸�
�*ng�c��SZۋg� M��0����{f���H�������2p�K���b�hz�TCX3`�;{2���Z�����ðlD�=��s��Z����7+o&6�I_	#;Y�kE���f33�rSQ�6DN.wpI�X�}@' z7�\����>���RT�k��z7��
5}� ޥ��y���Kv���)��[�<͢~]��r�� ^���M�x��._�)��:�Q����vhHb�g�Dy~��?:HD�s����p��V�gO�pB�A����Za$���2�s`!�P|�~l�W@���\d͘�zP��&�>0:�^��*�JB"�+�o]��!�<��-.'�Fl2��"32��N�y�v�πU�O��T��q F�u�W�Ҡ~���ޮ��[Y�/�\Z~;���G���h� \fpr��A����!�9m�`�xo��F�`s嘩5�2�[IM��:����)�wR^�>k��;���S��Hm-F���}eפc�i���O�> �T�m`��Z���N�_F�Um�/��Ȟ�إ!�y�Z��X���I�G��1��zl&���myP]es��n��gq�򠊼Q�Y׾��!4T����kȃd��l���(�]	�+P�M�h+a����lxk��<au�k��I��ʜl@[�lf�f�c�|�͑��`�n"P�O��<=��V��&X��zYorpT2cq����}}W�B������.��w�rZ��n:1'[�z+��k�����f�-!8��9�$���$�C.�|���$�*ѼE+s��h�̄Z�| K����n�O��tI�"#4�֛�5\�����Se��fS�����5:���Z�sI\���A? n?����l���I(��l�H'�9�Wr��_�% ��"�)�{��5� =c��?�(:����j|E�,���J��
��f�=�p��>6|�X��U���?��+Wxp��H��V�md�A��bmсt\�%�:6����/�8dv�}��F�:�g��ő��i���][�O��U�����Y��"���%�5��l��QT�ۤ�;e�.���f$�͠S������׿%@�����e�լTW�%���I+<
C1f5qݦ����j{J��,��vZ'��2�3v�˕�9�r�E��3e��HO���+,�,ڭ�6��H\똠d�ӌ��������B�ڭ8Z����vC�4��nQ* ��d�e�/𒚳��R�pxs��l�����|���o�Axv�I�Z�I 9>\�)���6��el3��Q�+Rz�������ǣN۠� �ѽ*�~Fu�I������f�R>� hP��F�6;F���W�!f��\���}1���);Ś�Fu��4����v���b{	�4�v?��)!+j�hȧC��i�����7�}������S�˘��z�ydI�b��(aW&c֯_]]�*�����&BߐcR+Y,?ۮ�k���ۓ\�\�0��Z�b���]=E9yld���?����h�� q��+��*��e�Pv�����t�+S"\�3�u���C5�YnG((T��ju�%d^`P�-����u���;wJ�{,�X�1S<D$Rv"��d��l�zq��+N��R�gExB.	�=��Ӧ�7�׆ϳ�o_�� t�T�]���#�ŗ+/�� �*��#�M��	(3/��c2��@u�n��	���1FJ�V���}�=}'�l�SҦ�2�N
���m���k1��;�Mۛ�\	���u9�nA��D_���$O������r�d���MI�!�:�X����?�Aq�P+k���4���u�I��j�BE�<w8`�AJ���8�7'��؋�+rE��h����H�q_.t���<��:���m��VK'0-�Yg���1���x1��7Ї�9�C�-�Q2�B��Q�p�%g���T͙l�N���`ۉaߙ�t��Br���{�E]��4����U��?!%Z��knp~s	���2ȡ�6�6��k�2S�>�P�+v��Y��a���ŽZ�*�#�=*�:s����.+������>`F4�Kdjɱ0D[�xX���/��5jo5��f=:��.�~��W'U��l"w+թ|55j�����;�����][a�y��/`c���_��2�Ɍ]��08�Nr0�^����'*َ�[�����c-�V�a�MDb�tC�N�wK5��6Jr���0Ld�g�����
�3uXJ�M�Q8��P���`��^�.șA�J'�+9�(�-U�<U�Ϊ����s��,�J�':W�đU Ot�}lɯL5 ��%2E$�,=aN���W�IL�d&C��̐n���&���rCrڄr-G:�yI`q�ٵ�#��v)-邈�9����s'"ь�Ǉ�AH�*�#Lcș��cm�~�w�&���^ tC 9$�?�������e����R�p	�T�&������J �r������}U\�<W�5�e�t}bb蠾 �{�X#�d���a��K�U�uZ�m�\��ה�I����܋�������.�������"�ڻ��XR	������%��4h�ᶰ��xpy���sl~�#^YJ�<r�.c[c�%�Lr��<Pdy��Xu�$T ���T�jD\��'xT�8�?����{u�?5��Je'�>Եq���ʴ�����26a��d:�p̙��5��v��pf�<$�����9�H���C�L��^�ǐX���T��R'��X��
��]Xʀ ��C�ZV���_b���T��J4�������/>�|��	���ٺ�;0�]	%�O���m�
��ʶl�T�̡E�F� �D�#��1Q���+�?���U�5�J�E'Q.M�Y�b	��R~%hJ�dҩB2,��>��֩�GP�� Z��X��ɿ,��7J�3^h��F���	���᷍'���Ј���t�Du�惲�C�L��
�X��)�=���9VXF>[�x�m/ѵ�^�@u�;���b��;DCo�r�sVI.�]�o8�_���%��=�Vui�zԵ�w�y1j9��!�H��ڥsGu�K�[|�w�e�j�����Q�8Q(?�}�ї1�C�s���|�=g�\���íB���OV��d�T� �<���o4�sUT oE9!C�m���B�"�z��.o6�j
@�J������KH�`5�j���yc����u7����3�/�fb
O8�Vwa���FŻz�&�k�h�kk�����ȃr�g2��(K��?����8E��z�>�Aj`��������he9h�^��=������T��7u)�/`��!5tSX��3|'� e�e�)V@!�x0�7���عV�!
K�4���MG�a�`��\�@����.BſzLٷfJ����x���ƍa)���d���i6z��B)�y�yڄG�&�Fn ?`[������D���c�2�̘cڞT�
m>M��4J��߂mK�JlCb�zл!������Wi͸K�7��Ɠ�q8�i)ѵp�f����l�O>8_,0>�f���K o�J��9��R��5E�n}�IV�+��ބPM�5H��*�)�璞�$� ��T�<ٗa��1�¾������L��H�p��o��}��Y�c洔 .Gb
�d;m��i�3�!�d�:|,$z��(K���_�3���%[���>Tkjxt���|���x�I���ur�-<uu����M���|m��޿_u\���?9�u�h�^�KԀm-Ǘ<��2&�g�ma<�,��L8��~�L�K8H���Hء��?�B���ZE'�7}�btKY�ŌȉNiEg�H���vBE�����A��?�@�ن�F�ݧR�b�C �����C�l;S%������x늦�J��*�rW�36���q)L{��"�b:���o����`�É]�楞��P���� C0��u h��P�)�o�C�)��:�<oMTSU/�n�~ɺ��4p�dV��Z�T��)���,�0^�/��݃���~uEËڤ>��!6�W�2��)�e��y�|��:a6��!�Z��*��
)?౭腐�F�~�i�-+b�{�M%��Zs�\��K�����t�%� ��
ct�s�j�k'D��x�e�c*y.e�33p��Eo{�G�����OR��$��;f��GY �5~<=�u��	�>��o���]otf.��b�S�nU�p���
���ܲ���X�\{Ai�d_�X���.��H=,[��噳�к�"�<�^|�]JW�4�b��i2F�#:�|�Ҥll�G�<�GӢ-ᖠ���x�&��N�w|���ٳ=ט̩���):�M�dL�5�#��SG�;���U����m�X��f����0;!�o��4�QJ���Q�u�S[���wr{*������
�w&J�3��_w�
m'������hLV&�[����;�P`�3e�؛:���l8�G)Ǣ�s��o}�fbH�a)�� �)��GKn�X��w�񬕴U����k�f�*׭c�WXh��|������́�P|�TR��В�W���ڂY��#4	��\~���cg7@h�)��b��{�JfcOa4e�����7�Yq�2�6��Ȋ�<ԏz#n�ՂqCۂ+PGC��>�>Z;��Id�1��c"�}��韞��~�%|d�D��]��5�������ؗ̊y>�7���/��`����8M��&�*�����`��&c+�Pc�|�*���cN8W}�~��ُ][E�&�E`O��-�<�s8��YqC��D�R3�Tэ0ȕ:ц�E������[�����H	�ķ�ɉX+E_؏�أ�¯�,=<Yϝ̜Dw�wXP0�2��5�=�݇ˎ�׾(ܘ���=�!��M(���f�հ���b����Z��;��r��<*/](���|� C�Ր�����h|�q\&,1����'iXvgv`��lU(���Zј��Cǔ�����5?�d�������.�C�/5mvLd�b{`����� �Lm�ήoH���f�lS�f[���V�>P[�y�w!_)�1��,�{�V�b��A��0�^����f)�dR���b[q~���]Ԟr��������)�Šn,��B�WÆ��,��4������\T�)A����~§ڲoC7�������0�I*�A��`�N�(p�������,l�P��a��?'��?D:W�a�D�Y 3� �X��`i���C�Qk��d��
�+����K���'�Y&�D1ٛu��z��b�O��Z�1Ys*�4Җҵ���X�����kmO�VC��N��WNV�����q!.�c�꼝]B�r�J zV_QkW��Q�,n��怮3
\�~�Æҍb�42���fp4ZO�t���d" $�٦�)�H�r\�Jz�=��c�%��D��8�g�jf̟*N%�B�2���Pǭ6$�7w�!ɍ��wT�=���HZv�2k7�_��VZ��b눘�p��Xf@ �y�zn��)���(=EO�ۦ!��5�yN���[��zF�����Fkۦ�A��)�o�������E��l{#>��}���E�,����7�i�ATol,Pu���e_D'���N[�������Q�1�;�#}<sJc�.�o$	��~�{�)�Ĕ=�N�?;7���ʝɎ�~���Ď	�i�*t[CQ#N�� �ɽW"n�f���S�6d������'%l-W Ȋ�y<�����7Ժn�(C�v��P���{� �����n�5M���J��[щ��H��f���\��0�J��C)����c$���G#�lj����x=�eI^��FV'b�$��6n\>2�Jт�Ӂ��l@�{2}�� ���6C�����a{jZ�E�R�?����]�Bֹ�@��2��ϖ���=�����1^��ꑤ�;���TA����5^$�˄����(�k�.�n]����
?�����2��Tʲd}�'��W@�;GZ����)��v�!&�Yv(S��z��4���&x��wIbН7<�H�lo���e��$yb��v�n3jT4����>ӊH��%�m?P4VVcU����F�$+٧�S�K1�~��S[i]��B+C��m�G�����-��&�ӫn^��fg��W����X~U�U�zbD�]�� Saj�N2����ۊ���>�d �7���H�~i���������Ǧ�:��g3�3]�c��P\)�[7��N�/�$V�c����Z�^�]6k�3^%��,D���*��������Ib�E��93+���D�~_RR������b��5�����	ž�>6�R�^v$���a>Ⱥ+�����r;9�&�	5=�,�����˭�1�����4e���G<G�
Y�D�,�Ia�A4��~qxbE�O��
���2�V��=�Sm\�ߎ���,�mR�;��˜aI��������''G�����2xZn�=�t��?-���fUj��q��3����Mk��ؕq{ E p�!n#�x_���֘��S��J��?�J:ߓX���,ø�/��s����	CQMKJH�3�e�S<�lgF�K[R$e��DIS5��W#�K�8KK�y�h=�ң.n�o�*z��54�[7C� �^� #�x�?Tw,�MF\ۄNcp�][��h�����@��d��r�l۫�m
��?�5�����I���
P��xA�oú9+V$�U[�!E���ǲ��OM�^� ��i푭%d;�ID-)y�KW�9C7�U�so�js!s;gƟ?���q���ڔ���ӊw4�J��\��߈�5n� d����Wl⹼K�iX��HR��4͉�\$��ˏ!�r�q�������"�;?����/�m��bo�)�WLb��Z<%C�I�WH?$�zp���E$���XJ3�=��(��1e�Z \\��ɔ޹ш@�Y�;MΠqX�B3!���Z�&�Y�h�5�3,��F '�����H�/+�bi�h��TYF��@�a����:w�a�j�6�x�ډz�ѓ� jP?�����³��:�yѢ�b�q�ge����u��k)i����A_�h�JA�{ ��#l^)�}�?9���O�(�z�nԑ(j��(� P�&�2"��9>��a�Ű�}+��@sޑ`�Щ�r��B}�{+l�����)�?�a���K�͛��T��������W��S�	�)��A���*������v������a���;gX�p�~����]��3��1��d����!(i��l��]P]�d�[_GӤ�-�\�jG��DE=�Wږ�9#1^퓙�!u��>��S�6ӏ-t1�K�4�y�P>��e��`b	ݱ�ٲ����!�k1,A����Y�І��ew̌��Y��奈�=۸Y4���nC����#�yI	!a��),g��so�w:꼿Z�&�i���d���D����kx/i�t�x��=C�q���w���?sz	WV�3q�cO�y���<;Y� �1��
3k�-�=�/�~QC-D�m�8�pI�Yl��媤r_t�zx�l��{+F�U�
��PE��oȿտ��Z��J�-�����'c�$� !�"v}��c~�03���I� %�<@��o��nՇUm���Qn�M-�	x	�����mS�g���d�X���^��XC��=&w���h��6t�׶�I�p�&���@K;�K��k��?��!�B>�JU�j�&���k͎�Z#�I�ϯ�z���́�I���^�۴��ٴ��6.��e�ԫ��.*���������B��ڑ���ڤ��������uǜ�����6MU��w� aѼwFڍ�+-ea#�O������B���k�`��3�\�}��3�)�[�>KR�z9�F~��o�,�P/�=���j�|�� m�EtE.�e���P��&����K9�>��OȊ?���w��}���3S݈NDe�{ƛ�7��w�*��R��+c�`sjf��M�����J����s�a1h!�g�0=��������Ot�#�=�́%�
G��d�{S7,��`�R0�/�(C���R�MF!�I�o��i�9|�@i���s��cXqv�C�^E ,�G�6ʶy��ᙘ����	nVFɡ��y��`8h�%EE�e��r,�1���$�nQ���7�?>A��X/�Wt,�6��zj�+��T�@,rA�\x9C��4�v�`��L%�y1��y��w�������}�����f>ځ�j�XY����mz�l	�K-��u����|��Mx��>��G���eEu�9S��d#�}-V�u�|�Vs��ai�-qE^0͒�CB{=Y���t}����;EwldC��;�N��k���}����b�,X��elY~Mo�M<�$��%�U��~=gB��
�؄�V#�	��	�B�5�M��q�i����&4��d�m�oz�]��Y��vQ��M��VyXR��#FH{|�Ac7��v�p9��e�̙Q�p�Ly�aY���r$��x/����hVz�!�y���2]�W�hm���.3�z�K��:=pV�2�ΰ�f�#]�c/ګ��`�zuH�l����S��Y;��_��A��M-2�c�h��,�0St��>Es��ZVX��M�������Rb62�9�O�#y�j8��"�)�WĽN�4��V�g����cXwm1�Jا0r|y�K��(�:�~ͱ�����y���:�M�ȩ��)��Ϳ���x:�ت�dߢm�"��*0�����/� 0NTqM�� 3�,�#� hQ2c���b(WEtSqT��r ��$2~�п�4�/��g���NŨ����� bT<�:�xb�t��C,i1�qkd�����ְ�P�ZIG��@}�%�8�� @���o�0�u[��:3rY�Vlut.�>»�v
�����#�`Ԛ��[{,�1�en�ق{��פ`����j�+s��>�f��9�wx
O/4W/��@��!�:(��V����#U��I�~1[F3A�K�����qR`�+��<V�t���R�V�������_2��|����������*���O�5@;��9�AW>�xQ������O�%�ό��
BJ�i_.�Q!���/��XR@?��n��?��Kq�7����-��F���cFh���)�gk�ҍ5���鑨A�O��՞R�42�c���.��8�w���?qf�����ḑ0�����.�&�I���J朲��N�� ]�	dT�0�8��
!z,%�0�ۍ(Q����R���Pr��b߸�yj�,�U  \��z�F��u��KZk��B�0t<jw�g*�m�9Yh�B�H�[�\(vΟ��Z��9��L���ԝJ@��и8�oYJM�
�9Ȃ7ۅ�-ې1�qE����MU������T;�#rr-^Ť�����]��O�L�#;*��PD
�$�[�����.�8ԕ��>�!��J�����S�CL�(�maI�ñ����jx"i��e#�M����L���N���)5�u|@h��=^��.]�aP�Gc��-6XӮn���#$�[�@G���*����s�<ip�W]���ثe��,F�/���$N��e���t~Ø�P����QO��F�;���JZ{=��0��Q92.��j4i���w��;�0S�CE�+��DZ���F#p	�n�<�0�o�)k�Y���?N���-���\խr�+�hkyQ"ي������7��>�)l++T��LV��D/��5$L��H�nӋ�!��a��J� �K��|a.�$�ٺ�K�Q��p�.}%��

�!Yy�N[,��2�Q���mt#Q��Yʏ>a�@m�m`vq��|=�KB{�-�a���T�g�0�<�4^|eC�Z�E�Ձґ�fD�4�)�V&0�ز�$���!�o�S�8B��%�kk��l;Q�� ����D��G6׏���RH���Ħ�j����7��3> �¥� ��C1�>���ӒDK��Z�(��Pi�r�6V��3f72u�u�yD����;ޙ�s��c^�����'�,s�)8����Ŋ@��W�'��<�ǽ�3L;\H�sCg�^x*&`�\�
L�k2R�T�7�q!$��q���8�le]Z{��8����E�;��9�ӨmH���
[�������3�w�r�a�<� ��ӹ��m�q31�	���#��7������	Ł�0h��j �Q��_�����/Rz�r�GK֪�w��[~�[�^�b ��-�@��mϜ�@<���FtP�\�g����U����Ő��bc�.�O�H�H�6F�ӕ�.�������0n�d��
�q)R�nh�J�C���LsSh�r������GUzK�Z���<I���
a}u���7%l
�5�^0|̣x�T���y$����P�����������	�n�4K�Y�:ʩ�&�\�(�t4M����'�κ'q<�T������!?�&Mhd9f����3���N�Б�|)�W	�P�K�,����UO��a���1U����5��w�"Xfux���A������QɎً�3�9d�#2�h!:E�X�9��Q�@�(�P�ɖ���3�ŪJ��bK���W��>�Qy�$��V����y��I:K�xq�4,���Z!>��DL\k0�h��k��K=( 	X,P�b���TL�#_��廙_��U$n+J_����л�/��H��6Z�I=�,����|��b�t�|�G|��ӡ����Q��y9Y��F�8`��"�P&)��TI�<�8��	�3���Ґ��)���1�47�H&�i���j�񉀩^�{s'��vPGI���?��6�x*r�pCF)ŕYlUyM@��A��B�����O�ɛ��R��;V�#������x�`�n��Ы���׭�5\w��^���Keȋ���>ܟ��v�L����ݚ���5�6��!>s��>1`N�씉����Q��
�?**����'������2�rl*|�󨔓q��~�t>:^>`�@2������${�r4j�A:|3��N*e7�~�'�.���7�a�1����������1;4�B`�	(��\	�H+��&�o�Â��Y�㉂i�?�Hw�L]\M\���,
���|�R�I�1����Q���.���}�5{*¿El���㮪X�2����7�f*��l��]ۇ�����͎ Z(�N�S]�&�݊d�Ϫ��L��#�3GdO�xiW�Pk��@��px�ʦ��SѮN?�fMy"�1��)ib���K���I%&���Ӳ܌
�F�D�����m/˼�f���<�fb��CX"�E����}_F�X�1��J�������:j�h���v���1�
*�fQ�\wǢ�hf����C�a)�Y��q�eI1;9J?���G?�>�Q��W��@�sA2ceУL�?(��AX|�����e������[�5r�|��C����H:tc����B�.I��:ɟ�e�7+�r|k���[�l l'�m�kԦnH��9I��ge���2�7q�|72�L��ׅ��E��<�3�$����RdH�_Se+�j�I�%F>��SF$�q�S��P�Z�D���t��|������Q�]`{���d<�ޠ��Yf�"�S6���ns�R���Ӹ6�I�خ�Ou$V�@�l��a�@�g��j\ko}�e���W]΁�6�I=��_d��:h nQ78x�Ţǜ�p�[]�����Ϻ��C%�${�}�?��u�+��1  1Hi��@hdsW/#�<c�>�L�o<��e�[P�ͭBZ@k�]�/�D��{Z���O5 �#Y��ݸ��jߌ혓��**��\a'���`2?���b�h��f2���%e��R^8�o_��#�O��O��ܷ�����ur�|Ĳ̇��]���kF������/�j�0?|kA�2�8�t[���6C����sݪ�r`<-�؞;븿�im����҃ꇊ�'_K*܎Lw^'b'88�I3O�M�@��5� �e������t<��ߞc�k&�B�~l�FhFB��N*�2��#ٖ�@R���w�9��]�W��U�A����!mEu+����^H��8��Z�\�d�� �a����������-*�M������Q�wr0�#��c�J�x<���W�ݐ�Y�b�f%m}���z�R�ȃ�*�ˬ�"7�?�����D*!����&5A|�Y��D�^�?Ԭ ����=b��h[�f#��QgK�cQ��M�N��u�CQ�]0JbP6-�#�6~-��e'ȹ��PI��`Tsp�5���#pV�9�L�!�⹓D|,����a���Q��C�J��yU*�/�G�ݻd��ZI
�&�Zڳ�N����qlX?[�"d��8���=ML�b��`�毽X�����$�tE�3�%�T���Jd��ΞLǟ���k:�}�zo�L%#���#��I;�x\Q^b( 3�_d��G�QP$v�����C��U��A��a�e�Ω`�|��cZ�Lޥ�����M�^R�K�	���4��
�����f���w������){��������J3cv�K=��Z��d���ox$�G{��.K���k[o#w��]/̧�N��s�0��xw��n��5*�����i�X1���(�=U)����PB��v�:[呀�V�qn�Ʋ���̂�R�`�4Kc4�	M��)rl8!�?��5�x�#�L�Z*OE�_�����0���9D�v��4��P�܀X�t�O�|*������L¶�w����-6��$��<�I6R��7��a;T��>L��T�^A�8��}F�t]UbA��������N��`(+<� {�9����L�u6#ǀ�%[Y&�?q���S"$Ϭ������ȴ��JJћ�]��*Ԩ���:ť�����R�!��搀�9cv�~S����&歾i�Zر�~k���/r��l��R��c�2}X���G����:L�8��v����#�_AA8�ةd��i���Dߤ�j��A�I�'b��H���zhs�8d�m�ͯ9���B��3[Cp�Pgu��tiK�T��t��
B@S ���!%Ӵi�_�;�8�.����)��r#��w���w;8e\�R�F������� �A����me�[eTs�/���7�.(6��3�ڻ6�����nx�����E6�(d����"w��G���Qq<�)�4h[�(�����̻1b�/�)����}���RJ�+ř7����!;E�
� l�&���$t�$���W5HC�|�V��*%W1C�Qe������_G�ږ^%>���^P��x���Y��Mj�~�"?M�o�rC���ۚ?8�/�]��ƛ�,�{���Vl5��F�2��kK�J�`=tS3�*]�t\�/�t��7���h��TȨX���v�[P�`+�V<Y��j%����;�閍o2W}@�I^�I��(����P߭*�%����B��ݢ#��՞�O�,�up� ��Z�y��I�V��]6��Ũ����-*�7�#_(�J��� o�+�釟�'(��v�4C�AW�V�v5����wH�j�F:.�,�"�6�Is�3�-�>�,�D<�&�0����'��x�!b �|��WV��?���8����b��7��J�G� ����LtW��[H��q����5nl�ߜ��\�OJ߽������.G�����/u��S�ª��B�}��!o)��!)�^�"*gm>���B	�	Sb�%��ch��0�U�3�:$>��V�*u�|d?�
�Ν�s�JS�O�H�m��Y�4w�#�d�w��6��
����P�"7��}h����]8�^���!y�f��@ķ���r]�I-	�9X<��lO�L�=�����%�1���)C�dzeWU�B�Y\��
�n��v��U�{�c��	����/"2�y=���<� &1�Ѡ�N<c��XB_�	�{�9 w�μ`1'�F�P�=̮�_���Dl�x?�crӴ��-�l�W���#zꅛ��������%5�+f�mY�+���n��8K��4�c�z�]"���[ �?(��r%��ܶ��+��k�_Iߜ|M^3Mc�ؽƼ��+��S��w�FZդ`0'����b*������֙Bwi�)?U��P��Y�D���F�Vr�yK���t_�6����eNa����6kMW���F��\��!��MJS��XQװ!~�}h�/�\�e��HeU����p���$|v/�~!�ei�z���0�d|Cb2��St�������ӝ5�"�$w��;��l�?����+���Zep�R�pL���`�¹W3£�TC��-��جv��x���੥��&r�#E v����Q�J�z-�,����p�������u� ���a�y��J��=�EւO!\r{(`���@σ���}�<�)p�L�ɷ�)�:]�A$
�.�+��λ�R���K6��K�a���R=�.�������1���ځ�5���[�ZA�.B`��
��煥�c{Z�mMǷ$��ł��biI�ȁ���U�]/lf8
P�7�������p�W���+}�YS��P�&}����L�Jt�HD`�SK�?��to�'w)U~�@����k��C-���]��p�ZKZ>@�%�g�lO��g��:l�A%���7�]�]�n?(2j��S���MN�Z#��V
Zi���ܒ�����z^�X��f?Zh���bnA���3���z��-��e����d5c�H��g_>��W���jQ5��"����砩Ο�/��G�[�G��u�ĸ��7S����?��,��X�������6�D$l����$ؔ]���1:��i��~b�k���N��H�4�A�X��X�u8�lH����Ɍ|����74Ze^�}'��L�잹�#S��I+ԗ0�=;I��.�8��6�6������h&���4F8t���LD6����,F��p��쿆�����~�j����"6�l��77�7�+�]Iq��J�T��t�`mm�؋!�{ķ�z��5@$����;���i*�<�t���S��̽xh8_KkRĻ���cm���>)$�#f��,���|� IW�@u��e���������rr�#��/�BkᘻJ>,A��2/}ln:!�V�؆�}��6�/�<�|&V^��s�XH-S[r��H#'jS���$�^�h�{���$1���hN6�D4X֥�t��LD�o(��O��W	�����(F]`���
D�q��e�+���P�s����+2W%O�����(w�ݙ�q:���Xp���dfj�|��v�~Q p���˨~���^U�a�T|ż��\w���t���#��g�����=��Nj{m݈����h�nG4z3��R٢?�5\���QS�>\C���A0�]ի��j��2�'�c�}?#<��V��)���Q��J� >L�S.*�+}�t��zi�8����r�<rn��E<ݍPo5M�U�H��/i��+r�� z��j�jw�A�k��8Arϝ�R��eˌ��Ѥ_T�z���j� jSʬ��)��/#�l

a����O{�]�2_Ne^���բd��[%�~����4{9�e�y
�/�[��
���7|������ƜAq�:J���H�ʦ��Z������3�_ O�!�_P��zr���o�Wr�0x�t�̔�F�qa��`����g�v�w5.I@�b&&T.�m��IĨ���jUX�*����[�c��#��85em�����AT�Ϳ(�CL����9Wc2�����[��r����[l'2}iOK�6&mC��1���.���h����(?��R]Cp�����A:#����/�㫟t!�d&�	OG��:9J���}=�O]	z�6c��9W]�^;� ��w4u�68�����F�����y�2	���+�q�g��lv��W�]{��t��K��u��@�V:AU9uA���o�31��� �|����K��ƀ_-�{~�W'z8�K�.��,�p sי��P�:m�F��T���&�:#۷ eG���azsl��ч8+���!�����;�� :��g�|j??�4����M@�]���=c�Mr�1���heh�$��$��L�m)z���U	��c�V(��O�mKy�S
%]��J0���Q!���x`�XtV,P5s�պ���X"�I�l�qN��]$��q/���ɁO*��	&�;��o~Gb�]�R�P���E}v��� /Lk���k>D#�y3d���\��G��VϮبE�i3&r�����]��
 ��z'�_��y?d�-b�-�\�4)�T��30M�K[	�(��Y0�ȡ�Ѷ��OSj��U ��D�&�nu��1�������_���+��c|x/駯W~�%�uX,��n���5+W���X��z
��f��V�'eGk�7� �K�Xo�:?�����?�+}�Qpv.l9��x)7î�]t�c�n��LW�f��
A�vÈV}��d�����<B'Q������SS�����h<1��pV��?#4
Mo�:ɿ��8�jສ�ؐ�CBSܺa&�[;�bԇ���]Hz@�68�'�IL!.?H_؜�Zm��s��f.�oo��i�<��~ɽ&�klE?V;���Q�zJ('PJ��"��������$^�tm
�A���(l[}\�����bJdYc-�Х��8�	��}�:���q�o!:w�����G�6
��Qp��Xe�$�-;���)�.��j�YH	�eT3�������9�jC̐O�Z����U� n�gx�q��_�_5��`J>���_��YL��P��k�#��kvm��F�9� ��lD�2� �?��.S��*^���C�(�5'(���#�OY3������"]=��>�ג��3��BWջx}L��Z�ƴ���jl��W-�	/�	��7gN'f��-pj�!8ሏih�j�|��.���A��b��d�k�b��nF�؅.L1�;�YG�4THDS�I�6U���؂z�]�H>�����m&��T}1��,��qi�^��seU����c�8��D�sI�uW6�Ğ�.�A���Ϫx�e�o#S��-]��h�0����iz,�ų��V�GR���߻�Bg�n��3,�GP�i{	��>@z�x����B��.���e�{��1��^H%*���
	8���)����_��}]���K��&W�w��Ao4f�e\E��K��!�#�:���&�� ��%��/ى|��B]N:I���HJ%s��I����G�}uj�q+H��&���~�j�zSd����gS�0�1�!��r?sa&ނ�d�/l�Űؑn��\�8c�t���ێ�غw˹n��|�&���|���w^M�b(5�{���5[C�ǨDn�[p}�Ꜳ)/�n�7�X9'd�gPE����_�#��3�z�R�|ysu�k�yTgv6�/D�}��k;|7[��=ğ��9ńj8@�gT�n�j]b���Ⱦ��ĥs�K��%���R��XA��$].�tZMb5�� ��q�[�ꎎ;�������^�~Ϲ��?�;	x].��Q������p�:�l���m[{,θ�5�����=3Ł����zl8.ϛN�g���ž��H��&�EƎx��s��m�u�dG�l�b�GW�\?"��_��e"�Baa�����c��	(r���%�IW�@�4�.�*`���mj�I)
�ri;`v��~|�C�{'3t��"C!~��*KEU���:O܌8ȭ�=�V�Y��� ,!�j��19*V
G���A}UD��(Mw%��/Kv�'.!�;*D���'�?FU����!��7� C�����6�:�mHD�����է(��bQ&g��Qc=��8�m���j1S�)���f�]�q��Wm 0&ZE�^��o*%��/�ı!�	(B�l���� NoeQ��B�C!����'��nU��=ZfQ���IC�&�K%�7���߭�ӳ"�k�59'0�l.~��T�ݩ\�e�Bʏ�,��r�>'���C+��f�@z��4N~U@
j�� tPTp����*����}��=sg��vd�w���ڬ�$�C���*Tv1ꋸ��/�|U\��r#pQ
���|^b�I���6@�׮H���Q��I�����Tp��-����*�[�cK�{Wu�=��1mq}�^�t���� �e�zd,�b�?^�����X���ߪ�����րH�G���`��s�z��`ՄA�wN �tl����R�:qr)��a�2ɧX� v}QJ���LX��Sp�����U�ͥ{�Pq�CT@�n3
�U��.�LÒ����̰�,�z���$y�%�D�c��(4��(1�kh�/�ҲR���[��WH,����%�7{�P��1�Qe�z���Ĉ��2nK��o�e�S�~�WM���o�|-؊70]����v �$�E�t����d�BdO�",W8<�S
�an�i���`�DJ"�&�U���&��(�V0y�>��{���S��)��{�8NQ�����:�cx[8��YX����iY��k?� 0\�gKfT�
��(ϐ�����5�`����r(H�vU_��G��K�\�0��y*Rq�$�MX���^@蕆�T%�<�Ik�0�����q�И/�,��
���sk���PS���l��Mw�L�vlXB��h[�A�����T%=�)� ��~�/�HR������3�R�Y�Z���
�u��.��Z��Ww*Q,�ދ��eTӪ%0�o|W\w��5�3.�
`��Uנ3��G
z|��)p�抉���ݐ��9�СWj�|bj&_�#/�D���k�aZ-��
b��ҡ���Hߢc�������ſ��V��g�[�Fh&)��Ŭ\uQU�_���LG��ݤ�Q��<�i}(�{#���kg1J���9ڼ�&�� e����/2LhZ�D��?k�6�^{�b3�Zw)j>��foT�7!&�Fxh��:�#�!+�Q@7���1>�"��-�_�Ԑ�K#TH��p]g%~�M����с�Zx��!�^��2 b�Y��RU-��'+@;�̨Q H��4�^���Op����o����/��)"��d���q�l5u����7�*�~�m��K@�SJku�Ack��^�����uv�|;�n�u1!�Oݿ�!r��BP��4P�r3A�~*wy�Q5S��-$@�T� A"崈5}�"�9|&�:h^�1�౔D��h��k"����9��M�>��|7A�
x7�eh2���D��β�`��Ǥ��Üҭ��Ͷ��%�?�tϟ����X���<������H))���}[�~B�Aƹ��d�*8'���(��K��U���G���ʀ�Ǽ�{ohhA��(��S��	�0J�b�):��]ɫ��Bo�6�ɢ��F�6���i8��o'W�ݨ��AP[��c��a�%cX%�)��G��eY��F����gb��#=u�$��ڧ���e�󮚁I�	!�#dK�t=����gҬ�`�T)t6�f(
���P�{D��p��DA�-�����{�����2��k�/�V0�����h��9�?C�e�
���,E���V�ce�#����HPvS���<HNXE�֊�����^nO���{Z�؝� ���͵�U9��7�Z�g0rU5��,��
�6�'YQH^jc�"Z��@]�V)a���x���	�f��Փ?�Hql�H��
�Q��Q�H�j� ��F��=T>�쵧L�3\�ܑ&�cH�����ky�'N/�S:�Ug⿱�E}H��y(�;��'�`��|�����~�h��*WZ�do$�,��u}�t������		�ښ������?^TR�$#Yo��6�g\����_����A?����t~Su;�x�u�����UI赂έ�z�5����5��V��y�A��;������i���G3/9�Y!b�FK	3�H2V�N�%s\��u�k��LL�nc|��s�C��X:k�Dr�8�^0��EĤh�0�.j�ɑ'��})��4�(��7���q�UZ����Vӱn?O��?_h1xO������B���n_4��4H�jE�=i,F�wx�y�p~oP�^���Й��	�X�M����k6$�H_�Z4����,���_@���9n}N���-ް�e=��-+^Ύ����ܺؑ�r��	R�z���<S�zs�.'�yf�Q���x�- �$h{��@��	������s�E>��E�
��U��sIT3�������$�p��m !��c��c�x�K�A������Y�aT:m�K�V�Fʑ������ML ��V���i�U���ob�T�&���<�k���z���o��W����U�����=���i�4־CDno��
�y���	��{CSڀT�ɏm#'���q�O���S�r�I���K��_H�`�#�D��#r��c6xE~bY�uXNB0H�B�ЖM�߈.2��r^�6)��3B'�u��Q�G6k��X_d�ɰ ��n�6�W���;�:��L$v5���e0�KJP=Dϕ燽�����q����Bx��ѳ�tC�|={�X;B�s�T4L�o�ͦ_ajv`��{eM���+"t��R�"��16��ޖc��K�(O��`���bd#�7N��S�%�(d��9x���ʴ���/Gj�௿RM�S�̳���c�/�H^�)�|��a���8�(J�����(���Rh�����jc���m�2�=ܱ��X[���Ax�9	{�jF`9�}"�%8��[��>.������+�@�����'��ð�۽e��w��ڰ,h]�7�O�P�Nd��t~O�(̓٥|�������Z��u.��-8EkY����+�'����ڤ�vj�Z��dO�4NZQm�G~�`��ı��"No�x�K�����$��Ua��m2�<�M�6/�+@�RC6�.��7)�ܱ�h�W"\GO�����n'�ȏ�]+%��<�TI>�*A�I����C.v΅����;�C
A�(��kX��hs�lq�R�����~Ҿ�zE0�.��i@�%�@�E�qp�)�|_8���%�e[ �����K����j�9��^m�M��M�J���Y��o,͝�䣊����8
[��K�� .:��,T1�Z��ie`y��
a�������a�Q� ���.���3�H�y���"�������p�i�wet��KX<h�\ �W�R�444kL���ѭ�V�B��D�N���Iড1Q����n5k��F(w@WT��)�[�=q�^a�
��c�@�-!��<6��}�lP�W�6��:]�6�W-<wh��{R�y:.�~9Lg�l���9C�Ym�a����ɠ;�XWSw_��K���rg=�jo%˳��a�8����)~�Oݯ�H�2׏�W��w�U�6�$�j�fJ�]e}��>&�GG�2Ŕ\*��G]��5��Qs4��i�3,�!�Q%�;o�5�y��+���@"(p
$.�õkg���n2AE�0�o�M�|\j�0��֧��]�a��bj�GA�iZc���HZ��A����9�Z�������O�nHz��r.�9�I��;(	�Ҽ��)�zP(t㟍��D�����׬Y�c����-�8��E��q����	�&�)��m/,f"�i�4���N%��ze�q�9��n��@�1���ޗjR�T̡3�/ȫ1>�r�]:�;6'^yO����bc�YL��#�/���F�F-��f]8����:�}W���q#"<�Bdǻ�=� u\#R�S?�����)3�#n���+�Fy멵>��pZo��u7poG�}x*.r�/I%-�"�(�UԳB��'�,G:Q��H��͑��Y�a��-̝۪y���PW|g�'�P�\�e������e�imn|k�$�#ŝ3Y�T���Q�ŁM����Ʈ�i8T�JT����rT����\n"��zò�'�D���=�0��܇�R��0�{ΚT�U=��]�a�>!#�U����9`���r/�Ĥ���,��2e��[{��y�Xf�~�z@8Y5�B������m�h���D�<Ϳ�QS���y���Tp����s��F��T �
�u�i� �݅3��,~���O��Ą봧p�Y�ᦄ����5~65F*���I�������5J�@$	_RǚFg1";��3A�m��p��S �O~%Gͧ�T�k�v1y"��2u�-��t����� @���$�oJ�rwa�����T����W֮�'lZ�Μ�hA�=�y�Q����}1�{����m��c��!��Š�]�O\�����炚�OL�[ ����g7�	Q�=a(�����_��C�P�b���݌��p�e�2�y��� ���
͠�h��k��UJD��U�Fg�[$�ϋ�wڤ}��2)RJ���ѱ�+~b�d��� ��Kq�7� �hQw�J<��ʽv�)x����_w;鞕HD�8c�[�í�I�n�6X���O ��N�Nk�}�'��o7s��gJ�d�����j*?��nzd��@.[殹�hiͧA�znA{C�M��B
=ԅ[ύ��a������"�&���aR|*�=�-ŭ6��x]6k)����0�
��聦��l�@�2�⚱i�5h��C}�B�<��1�7� �R�#���r�T�eK�*m����cK�^��fkm�4����	0�]�����FezVЏ�K�Kh���2��wTZY��Pb!�Z��6��m���^:�H��KPl�f��rB�G��&�����QW�yv�JW�T0�\������I'In���ک���>~�z�x�JD� �Qh�-O�����	(@��N旊���ű�6Y��^�ֽ�9SB�$�#&��F�젣)ERzOj	;T?�w���i]7���@-6��󕹒 ��I«@ԇ�D�h^���@�@@6�p�i	u�K����ۚ���
�\Pa�c��^Yg�f(�6��s8	�Ǒ�Q@���5������ṅ�f���<�h� W\'���i4%Y���e�t���2f_u-�Τq���YXb����ö�;�֗�ı��d�z��p�De�B�J:��f�OE����-�&��%l�j&U�`A���㾇���ܕj�pn��hB�|ߍE<�3������+���G-�²2��վ#�
��T�g�z����֧ɳ� t+Hx���>���|�ϰ��X#�!j_ʀu:cÔ�Ե���D`�#�����+e7�m�E�c��Q�S�$n���@U�[h�|�T.�3ӟ���3P8z��>��xk��������-&�"�|D7��5�/����
�|/y�:��F^��=�|�=��T�-ގ���󸺉q�����ʈ�q�G��ҧWײS%��/Qe�6�J��(%���������1F+���2B��
�A�pŽƵ'��ކ'P��[0[��f��/�b�j���Ջ��+r7-�Hǆu���+��KCeIwR�8��aX '�Y���J<Z���#&:l1m�#�LՕ�ct3��R�X��H�������͊�2�t4}��Y*ٞ���D�w=�q{�\;���N�[�����x��T`�c�K��#y�L�����6N�	�{&֎,�� �j�S�����J�X�Fr�9��	D�)�H�"�� �����u�4�i���h���V�ަJ6�(�a�j����:�	.u��	*�����-C���!Y�]� �<��
�O���D6���#sx��:;�w�3W�S��3+s�[�*m��8���D�~4e���:rX�qX(��^�N֕��"o5�<5e�)é�R��F;�5�� �	H1=|�E~��B���~�On���Lqxč��[P��������e#����Co4Z$�"��M���_5<u�ٚ�djK�FgY�P��'�9��Y."��n_��uKo�b����4�t;>�H����1vW˧4qi2�`iS��9���gG�Pб)Ih�=A�l�<b����i�ua��I��=�4��
k�>����_����"'#��N9�+�m�l�l)���N2�'M�a�k/�c�#�:�Ǹ�����r���ԗn��v5<���t~01(H��=��������A�[��;qM��?j�4�i�9Aj�w�
r�W�e<?~�o��KJX0�	e���^������MK#�
�:W�"�:��<_`5�d�L8vɲ�ن82��e�͟m��'FP$��ӎjD�X�~$kЎ�?�Ƌ� �7�~�=���_Ed5�b��L����_Tf�v�`�=�+7{9Qu���;1���:j�򑄉��6/����0�pK���2��mw|F�9�n�%���b�e���p/�H�z�us��+�Sj�a -��Uz!`�EJ"��Q�Ɉp��'	��@�;�1&��Wr��{�����w�������A��I�4��p�@)�U�+�C�[D+��X~�:sRH.��q�o��ѷ�q��s)X(g�q��a3��U�ĀQ�I!�n�؜g�A�N�ǳD�$���h��	"r��ҹGZbw�L!�xY]��Gz��6
��8�z�Jo~G.A��фB�C���~��.W�F��,v����T}�V!���W�����/2�m�KܹJ�`M��gf���&	^_?Z=��:�d�o�Y"!=t������\ǰ��1�Z��<)�5�z�hCSW��&T�$�*�&j1)H�0I�{�}���( ��Q���B�K��<־t�f ì�x4I����4�YZu���M��ѪL�;�C;qIи�,���_�p!s�I;����g�%<�ƽ�j���H2�P��XU�:)Dp�sw��	�{���τ|>�w��/���O�н��Ó��o�i�T~ojaȧ�����x@|���M ��(Dd���%i>�  � W��G��[�@�]�Na��v[���p��Fl~�r�� K�כ�,�er�����7��ΎA��K)��`G�� $ W��%�]ݽx�@n�e�	g����k�cO�tΛ{�+�5�'	>T·��b\�{��ѽf��=�߫f}~�.�̖����v��Rr5���y��%�[�fu��L�tq��H��p?�VO��E2��x�	]��$��]�M�p����?�,&#�%`04$en�n>�,�'u�W�U��llN�Ny�.$U�o^7�a9s5Lں�3�s=�3�|C���H ς���`ER�T�� �hO%��l��ȧ��쮛h�:���7U���P�nu���N�V|G��/m
��F�����L�T@%�cv��_3�5c�,"��!��^Q H�Lǳ�N���Dp��I�U-pve)�-�y?�ڞHA��7�+��g�R���b&���� I�5�d�w�N.�<����"���+�r�,a�L�O��O餕����9�`v�0b��^�^QTTˆ���I-����gV�8�
�Q��5�Fc"q1�AѦ4�2�*n��l�Y4��tf��W��K���N̚�"[; ���lЮ�y~�?�U(��a<@a���!oG��`�TrQ*Cٽi�j�p�l���ï���Tege"�����r/]�ϗ���E���ב7��OE�#����;��;�W�?�{̯[�`Ml�5�u���?b���e�2Aْ4��?��j/s�Z곽T2ȕ�]&!?�~$��a8P��R[���c����hG�X�C�6�G�Eu�	2�u�C�S���f���KKl�������Y�Vof�Y��r�,	h��b�u���q� y��|��&M^�2!U�f;��:hn���T06x�JɈ_i��cԷ'�g)���Hۈ=���sU�wx+�,�i8�T�5EU��~Qx<HD��@O�ʯs�4��ڔ���� �N+���w~�<����~��%x����6N� ĄP��/��=?oTCϮ{Fjf)�U�L:���V����o˼��^ڛ��2aS��J���>�0=N��[w��� Ń�]���Y?>r���\�m�!<�Rb����>i�Ϣ�䮙�Q��k��n���_Xq�Ih8d.�q��ۢ���_�9ś<̍���۽PI]o���4���ė	P�����6����A�$����O�}�u� C)������=�Pm""��Z^�[r��ꂕ-{�@�������ܼ���c-E;k(����ݢ�=����p��r���7�X��r�k�x�t�Ϟ$&���l
���#Ѹ�0�
��}/G����qG���ɟa<�z�(� 5�����[TVRԞ|A����}�S�����#tn�â��m�I�])3���XV�#3�tM8|�Z9!�6�l�o��w E���7�k�#������˳�������h9k���'ˋ��H�2,@�������8۱�k&�O�n}/��c땗х	�B=�M������ 9��R
|�A|S�`]P�Տ���_��t�S?���1�ݵy��r��j�-Ҫ��߱������r�����5EU�k�~��ۓ�"�O|OM�v�G�~�
t�sQ�A�)[ԥ���W�-�x�^�퇘�l�=�W�Qk��,��Nxe���<��3�j��H�$���s���\��,�rw��%��r��e�|��˪GQ�ŠWj<R��@͜��5�z7C�y a��cf���U*lƟ(�5���Ό��{7�6[��2�\�G��0p��D��&8���4���ń��>
�nv�9�w��I�td<ބP�5u����h{[��3���i� o�g�a�*��ٸ������	��r�^��~��Z�҂\��^������O
)�<����v���E �p�E5����I���i2G�����S�ٮc#P㭾�����^>�@��@U�И���6�rνT'Hd�k�뷡]A���%����A=u��K ��#cju$�U.3�Ր/��� �V��§�m�<S<��Ū�aI&�]l2�,�����|�ZM%ʯTcB�^�8�R�J6��+�#Z3"�!��۠�t:�'�H��z"������Gh ��$�y��e8j�C�����dD>��'V�T���͋���7Vdt����W='$Z8V��_7QatFȱV��������׶�oL�iJ&-����[х�q����l����gd��б��[�"Q�{������Gݹ�\> �8W����
�Et�z���K��I�"fx����Gb~3��^��ܠ����!Eq�l�l�S};T&'(����$�/�şTE��o5������?�(�RFG�,�A��.7�0	Y҆ŀ�	��Y�>�k3�{��5��|�;�d�?bi�k�Un���^4"u�s�35�
��eI��-����N��b)U�rgu�A�.��x�L�c���@�5KX��<�a~�Ig9�{�;].V�v��*X��%w!*�]z�4��M(���6#���~'V$�����~ �%ː�"�����G�ͷ}�I�#U���D#����>�I�]�8�L��o��d�
7Ρ�s3���F���'����L<#��a�p���J����'�r��R1[趄%6���w2Y�6�⇑��V����k�#���yŅg�@Є�`���Ui$R;�)�I
��щ�국	��R#��������F�t�g���,9�;D��QI������KgO��7�O�A��5_��0oe��J�/V��G����٫',h+t��u�m2��,�4�D�T�|75�uD�K,4�7I���R���ӧ�R��}�AI���z�I�g	횥�X�j����0"F�ߡ�̸U٩n������#G�X�u ��{���kB�77f���|A U*q���xl7rj,��E�7������c�ƮX"�F�E�7��b_�zC0Ԉ u��ۖ��lF7���	+/���[��ۛ�������|I��;���J0M��N��@�G�0gС?��#0�wJa�	�@�"ZL�%4�m"��g��K6�(D?�|Y�W< 8�LM-"k?�o�,
����jQ�ճ��R����W�M^ ��6��t6+|%��c�S2�׃�U.׾������.^x�����$�Q,N���d���D���aGc1~0��h*��b�r�J��!i^��[��"�+nz����V!\s�-�f��3�8H���[<�6~�(avx�]�CY�o\j�!T���Ey�{d�/�KP�� �� X,"�ړ��{e�ڲ���$�$#fS�Ϡ�N#��:�X�d|�i�9����-��{���֒K� �@$&!�|miXg;��`u��bR�=�J����v�iN��눓�q���*��+�5��4)!C�>�j���p��زG��<\����є�x{ϚЂ�'����wy,8����Rw���#A(���S�kd+�	+��+v뱸����x������*`BJYE�Zx��>�G&s(��f`DE�5�S����]��x�M�e@'��UK"v�ťu��^K�16�ɗ,mU�V$�4�8����/��n�`�I}m;а��;Iz��H2�z�Ǘ�~�8��-���U����ްu[�vʃX��K~k8&A�� �����ѡ
�i���$������.���ͪOT�@Bs���t�̌���q�S�j�x���p�i`2w@+���X�+#^�!���h���H��[�9��Őm;ؓ<{騞����#�(f�jo�*��� ���A�ן���^ѳ�[�I�` d���e������S����L�ߺm�<{)�"F���^�a�������
����n�A��.��,�3�?����փ�3�mQ��1+{�M�RUyk:i�Nz"s�J�s
A�3u�T�G@O��x�c�ov
C��e8�{!S�����۝s�Y6Z@6_gf��
_?�"�>m�\�4��?���������S�W���s�E�ڢ��x�t�4n�Xۘ{��v�G�(k;#��!o����^]%�HNY\���=y�S�"�_��V�@� d4��N�y8ߣ��&�|JPJdS�fvo�2ר�;���x���n�KZ}m�DE���e�7�g�A�c�Pa�bq�nL�!���ޅ������ӳ� �,�h���*g��WѤ�	��ҫ����b�����뙏���i�3�0�Xht���RFo�4E����TDu1�Ĥ��K�zF�3S��=ȧH�#�f8��/��t�6h,''#�U��c�<��Q���N���F4(�34���RͲ\;Y�����b��ޯ���"I�ѓ�$�'�I�6��0��!�\�ʍ��j�`��Lgh����f�l|���y�ʑ�8��8q�v����$Sl��Jпm}̏l�z�����uI
i}֤n����C���GH��P*.�y��.�5��خ+2uڭC����Yu'��2�}7�E�|ZD��8z�d3��e=#�S���>���d���Z�%����C���C� � 5*���BC+L����z�	C|l �`{&]>�_FmV/gy�}��y�n@q0"���j��c����!�]�@c��BuY�S��o�d�e�_Kw��H��	�E������aUT\�-7d ���[�k�8M�"C�_n[F�E�^q狼&�Y�pp`����Sc��[-\�Q�rF�H��aq�v{�
M�Q]rcvjYˇJ��0 |��9j舴���������t>�D�gqZ8w-����JA���B�����a��0��6wq���AQ`���FW��T�����F��� ����pE�2�ͷH�Mb���$��/�&���h�%��McSK����9�io��}ï�1VES�ӣ����#�������벹�X�ŜNK?�s#�K�c#g�p`�
���s�5*���2ːW���qB����Έ�0���nt~�ݔ�;o��9�&@	=��eGp�%�L��t��4..�e���6qN�C�Rr#�N��܀�)Җ�"���x|�fE"�'h7�� l3�χ���,��d�_7V��6s��s����o�M��.�h$��S���f";������d��I�s����Qo\~�p!a�E�����W���f\�y)���	RoBm�ȹ���Ho\�o�3�@c�B���)��I�4�/���� XA�
Ǝ_�K�w�kN��g�N-m�i�q.�~{�U�2����%��);8��"K	;d�����h��K?�2�'W��62��>�o ��*F�i�N\+L��O�3f���L��K�s��2~�Sڞ#���q��iX�~qhE����k���y��]���Wl^J���]H�|9C9{�t���gm�ӛK�?��Wr�Y�oϸIiw�fMJ�;�j��n��h�D>��}�E'B"�����`� �BeP=�j���(��;Η�F��1�竡?�褖 �y��cT�uWCω}������ӷc��:�Gh�Ǿ�*V���On5ǅ��8�0I>�w�5�Vn7"3Xչ����x�<�#���Αs��F�"S�]S�ćg\��Dm�a�l�{�j���k�H�8=8kS���F�\"�m�bW��4�p�"c���a0ӲNP�Ik\��~�7�U?J9ђ�V��n.x��ZU�^u�OT�+�7��4Fr�P�J�[_H�߾�,!3o�+�u 9��G7]Z�g����K��V_�,?��f��&�ܥ�~�9��è��}Ey��W���[A��Ћ��.	����4���G��ݑOo��ꯉ8|�����ު!@JF��B��2瑡[k�4�Q��`��2�����7�o��!���7�<�1"���0K�7nn)s|<����$��wcH�,� ��[�WG	�(��|!��c�����?����r"49bϾ$J��d
�-1"Lʌ��()��	��r)7�-���1`�n�ßK�~3�\`��S[b
Gr���a�#mSL���|�Ei���?q� h5?�פǎ�\��D�܂� �`B�>%Hs��0aK9�����1a� :�6t�v����^���U��fҺJ2�G�kX�dP��b�o�����������N���𘳩��nT�y=����CQ�	V�jzUyT_���ր��Jӛ��'��%^'�'�X�Ѣ#% ��K�	��J![@�.K��d7�\�ge�Fݳ��a���5��I ��֓p��s�FNɪ�I���B�Vέ��>ώ9��u>{U�VEǲ�p����8�v��ڒ�@'�B�� �ު����P��ΐH!ծҭW��I��{�:���C4�(W����,�3%�oy��뿬����Oy�����M�� :��[�v���j��o�_���Fר@��ӻ��}H�[P�FaQAFϺ�|c�zZ��ϖ� ��,S�7ƌ���ed8�%-_��
�R*g��:�A��o�FB����'����5��>9	�5�暂���W�pGk�����7�ň9��^e.�ZR����:'�m��6�vy��CE9�#F	E�Z��I) �z��=����ps�'4ؖb����=����n�؞��Fc%��ʊ���[]h�=����$"y�F�'���;���E���&�������H�o�zIX�Ԗ[�)��7�CLT_��=3!�e���"_�E���x�I�%�/8RF��$z!�� ֞w�' l+Na�f{�YhbFj@;�md\"�Ɛ���)�	�#p��+Q3:�#��"l]��6$k�X�DkP��"�xX�T}8(��q�kB��������+8�FK��P�&/|z���j꣤g0@��n��b/��~�C;Hr�4s���V�i������U��˺�z�Ή��q<�G���l���{b�@Ա(*6�4�Lf	��b*�f�
²{=q%���)��IL�L\e�1�;fc�k.��M>�",�F՛���Z��I"MA�o��w<�;F�f���d���,4��X�`��5Q�iT3͸�[fV�m,vJxC���G8��q����}pY#��#�\�ը�����e�b�n�P,C�嫔�/$�����*`mC@䤺��9�B�b��cO��@��;������mm�S����ظ��T�p���,)C�*�w�u�k/�a`-��(��2Q�5��#�16���\��]&�2��۟3��p������Fۈ�����z�k�n��+i&r������&Cp�>ҩt��ʰ�WI�D���c���.��]���6����Ca?�����6�����Վ�=P1�97P�p�tF���������}Mt_�YI�w0��x�}Ȩ+��1 j���"��|bppӟN*���+R����,�qn��%�  HU�,��?-����V���Kv�fϚ���{�8#V���_	��� ����(�E�9���13]����q���aG��q��U�H�u�#���򱜁�q��x��&UkSw�ʑ�Px~U�� � :q�HE`~��I��z���y4���d�� s�å�}�Q�rhp���~Q�C����>����).�����A���a�} �B,s9^A�1�v��Y]��(�$ߡ!ڊ�R��TM�n\|����:_b�d��I��J�� ��� ��-�\k�]��i���F���-��Ac�n�U.j�� x��ɂ=���a�8.�Ȅ�!�B��E!&�d#.$������'�� �2�;VK���K�����Xu,g�{�Ͳ�V��q�T����pxW��qϑ��=i�79B
�-gP��w�6�zӄ`��0�^7͍Bڋ�7%�h\lM��&�y�p(�R\����!'D��������=r��o�f��؆��LPi�	��8	��z��g���T����z�5i#x>�D[���Ca�1[(��F[g]3G�艽;SʇX����\�ٮF[[�"��s)�2'���U�yH��FJ�7���Ġ��	s���Q��"?~lղt���O��1[4���%�승w�1r/ԇnJ���i��%�9<��35Q\}n
�j:H��`F���z�
*!ى5�.�y��yb{ｿw��VCN�����[��f���IC��+em��?��?K��W�q> TA>!L��	����,{6�lx���y�;��yz��^�֭���:g�x�$�p$y,�_����&p�T|�ӑq�U1(<-��Ϋ�<ܚ��X�`8 �69��Q�b�����_x�2|ռhd�(�\jz@�X��>�d�k�[�%��8u���T�H�t�\VQܸI���g'�:2]gNu�� ���G.�-�ik2�6U]��4��*�t
W#�����#��M�Lj�d/{��bt¯�)Y����
F�,���bT4��x�󉅼k۟j��D6>�g.gO���2���<�����._�0_�̗���$x��G�-}5�Kk�C��̦0�����?���N¦�k�]����u!�_�eXwza�Cw�O�`O�|���I�792�FQ�o�i!�G��}�)����gs3C�O�L���a$E�V2�I�,l�o��&FY��j��r��/"��d>�w%��q��f9��mkwa=T���o���S=�#y��(![)�r�i�����9zu����\�O>�Y^m��P�zJ��|����*T�H�2���`��@W�	� 
�Ѯ(.�[�S�tl��uB��֪�H9N�ʴy�R�H�h�=_�H���v�7pA��'�ݗc�nI6�c�j������ӷ�_<*59w�<]��8����ĭ��=�5^v>���.�G�1�Zn�o��I���7�'�9�S�?�$����$H<� 0�ޞ�+vzB��,J6<i~�VAF��u\oK3�tm�	��9��vْ:���������O\�u�s�,
y����,K���1?+�	 Sv������?��f�d��<��R5b�ߜ�Tc�~$��ub�I~@ E.+�����j[_����(��Ν3�|<��_"ԇ�e��@%��p�L��y���7#�_(|���T��Va�O�������Bug˗鷙5�-�����hS��N�
�S<#{�[+m���8�t�%'
�q�w'8m����gKR'�F\PU�'�,.�:�[B����Eb�
�#,�e��Z�w��3� ����'[4ohÆ �K�k�E��_��+?n�z��}��A-Q[=�u���̞���� ����D�Hu����_J �f+��*� ���Z�n#���=s����{��?�{qmR��d��4��۵Ɯ�P�<��j����d�Np��w ��nd����wUU�k��&uti��ݶc�[��`pk��S��N=b7��O��m��I֛nV���A "#�������c��4Q���BO@��m���p���D�@�Jv���2r#��5"���9�Z]G���o̫�n;_� lu� ΠM�=�I���A_�;�>P��l�w]����FGF�|�`S�*�<��xL�YexI�if"�OYQ�G���q��}��#��G���G�=�'�����;ݘ3��}	t��ɩ��¶���8���j��l.�+/�,-�_��|)��}w���;>eF�a�N�5��7�٥Q}`��V���~H}\>����k������s��v�ﰴ�O#ꚩv4Iɬ���[b�]I�)foJ���*�^���4+ j웝j1qҸ��vV�y�e�S�[M&��e�B�?= �#�3O0�ۚDUNr_��\��1���H����Ì��b�C1p���de��&P���� )O�8�LM�i�fo�[cH�4�=�*Z�7���H�3�<+^��w��r��HM&~�5�`�B���Y#��8����"���<]s`�3�N&O��o�,�P�3`��" �W�ϳPkNk�laH��7fs�f�=F ϒ��k���8?`S������B�׉�k��eW��h��!��Phkz	Y�o�?hv��<d������^�7��*���7&��6���t��0��
�6�ٚ�h�#X0H�2��֐�Bh%$=`�<%uj������ų�I��������-��A-r��1�MC$<����N ���_�5�$|�'SL+��Ykmx��xı��s�^u�S����ס��/�B�N�ZF�b�g�����j�_q���=&�%��Y5�"�5h�2��c@`^Q1�u�8�/S���r��~��V�M�Ւ���Z.Zv�g������pD+���|�z�rOӢ�1i�%ZgT��"Z��jtx�K69sG ��s��1��[.��C�!Й��S80��Bw�u� ီΪTF/;���iʄ!���^��@9X	�f��͓��)��Wr�6��!���TVi}cw�]:���ψ�Ҭ�ݻ��f�Y�Ȝտ^�H!!Jn��@y"��������%�,���j��4"a�it+���E^L�|¥�KyC�?Jp�ۥh3=m�BNdR�����Ķ�G�������Ӟ���\�xty'��_���ּ�V���^��������Zl�kj��&�� E�rw�Ѝ������<�< np�����qQ���p>q2�E��"�3����#X�p�AR0YR��Oj ��F�7��4�%y�T�Ӕ����	|4�?

d�%Rv2�2n5`��*.�T˖�R˵��5u�\�Hu]U���Y'�d�xJ�yה]�5.�"N�׫��XI*PRT��q׺� �9-�{Os$�+���Ǻ�*R9���IL�>;S��+�o���3o��l���N������^$~ϰ�n���!�������D(b���\�J|N�����t;�\ĺ��n#�l�E���!a�4��Lf�ЗOO'�͏�9`=�;�̷p��B螹PqXf�i;�e&�B�_���SNg�au�_��?mYur��I�/ �">�nXK�ro�0��}�	�#�Ħ�&1�pĂL�V�@�Z��oY�LO_�O=����V�j�J�h��(Z7�BgZ�y MoM��B,4�j��$)�SR4�F����N0:'~Sh�,L��&���d�H�S@�y�z>2��ȗ7n�n�����k��}M�~��RWy��;e�./�.䳘D�fK���o�m�H�Cd%E�g9wQG#�Ԉ���]�(��4)q��~w����?#�U0_��� z��Z)Ԡ�Qd#C���ڮ?���|Eŉ��e�t���6�S� ��#� �F؎
J�w%E3��ե�@Šd��$�_���^2%٢��v3�STK7���W�� .zϾ�hg.h�jt�٭���ϕ�����
�m������;{�}����87˂�)~!k��4%'K��)q>:.�=��1��1�S��S)�?��?�Qld�Ӳ���i?�G���C8���IN��Ͳp5�$�g���P�c�m�����B�]@�7�S��MAnbt��\�߀�?��Rn���gg��K_ɶF��*�Nv�����
�j��r�٭�⌧'2�q=ad����ǌ	�S#߉�j��r��|&�[
�����a�`yƌ�~��a~���|���M���ˉ��x�{�]:��.M֟�{��~�&�M��>���"�J���,��x��!7^��%�N4�8�3a�Nu@�(9�t�zC&& SpppG��!ڳA���K��ש�>�&	u��(�W�l�j��T����*��Kg�E/�-��gD�\���6E"4�c�H������]�(���1����BUJ��_1J�q���P��	���iQ�FsS7�S'U��V�<��yƢ��:�8k���=e���+!�OٱMi&X2���=�"3��s$j�K�	�?U�g�y}ܻ8^Z��S�`*iq��"	"\kj^�D��߲M��s�������?xL��\C�����|3F�w�b��O������V���"�,���ZV�tФY��[l����dd�r���W���\�����m£�D<a����2�h��Z������~U*����i�ϋ(��ʕ�G?/�
�%���0m���r���}L9�Ǖ�������u�����=��=��l��6^Q���͈��l��6'�� ���<v��3`gO����p�"��)	�,�/��撌�<i�����6s�1x�?f����(:�������r�|�?���q�G��9��a�*���8�`�lȐ�:�L<����$}yU�S��w��
��R	2��3�.\�9��h�������;㚾��q����o�q�l��s��G�y���jR˲b�.x�2�2� v��/t��5;��O}��`jh�Q͐Q˓(�-���#�
T���H~���A�:ž}�>��ގ��$��*>���0Ұi[+�U(ä�z�J&[�s��/�%9��C��r�8����x�BV,�f���<��7�z�ڈ]Ő��B�{��`�J�x"��y@�:��S$g�\<��v��V�V�W
�4hVm��_&�W���(�'m��+*�Y}l;�Sџ�۴A�J�X�X���/@zl��XuM^�pJ�o��\�{!?Q�4������Hl�p�(����i���z��;�e-���mg�ך���{J�B�
 B��NO8L���_�a�OW{O�4�Ǩ"w�S���$���5rD��+C�2��m���J���X^��H��f��"�_�q�3�؞��j��s��U*#�L�k�V�DĚ���^����.jY�*�JyM��P9���UY-����r�� 8�;��v^)�#A�Z�r��!Пiu�agE��d�&vQ���e�kx�U���s�����!7%����>����8,����]v��8|YNJ���h6Sg�x���[צt�#s{mpc�N'SS��g˅y�� 4���Ñ�'�?��Վ�Zb�Q���J/5�������4�-e:��	)*���3TRb�-��v��]BR���W���\����q^�k�����g-f}Yٵ��1����n"ס8 ,׽!#�qDl�BxBB�}��P����KÇ�"�Z���M�e�Q[�+�$lҁ\�":�=����)�%��ǕX
��]�Κ��-����7i!Y�=����������Fv��N˿붔���j�� `�UV������*{2&���%Ǿ�� ���8����5���{�5��cJ�8��N���Q�����5#��d���Uma�@N�2�*-���(��A>��(��R?��ڭv�ޥ�� ���:��kh<��~=}�����2_���PG��A���Ӕ��z���p�v;d(Z�V?}�n!��Ĺ�����es�ʨM�~�ǐ�>��g�V�yӇLo��ˌ_@�꒣X��D"�[b�?��.G�O0ƋdTd��}�-vp����?�X,�X��"<�������H
F��%���"�?�
wS�#-�n�	*$چ�� M��N,Pz�v�cg8͐��FH~�� �Ԑ1 <����By�*���(���
��6�y|oR�7E�5]z�44�����C�DT,��P��m�.����T�Yob�b�yk�5:7&U�+�yb���3��U|�2"�}���b�����iq���v��g���Ӥ��t��d��T�`���B)�OB|��z��t�
"p�(z�����[��CsP��T���	j��;UW߮&�Y�������c�ˑ;�n����D�8��N��|���&��ư��*L�|�2��{;+���D���Rh�O��t�!x��ĖL��������e��� ���L ����o��3g�x+�'��A�(^�\ B䟩�(�����)�hd&{,�=��R��uiB���iL`<�,uc�=s�Nݯ</�$��5��բQ1�=$+ϑ�~�)�+��f-�<�F"ՠY���j�8'p����Y��4�N��d$xMs��#=dŲ��;=��)T$���ӳFe$���u^t
Rs��L�{1]lO]h���E�n�vֺV�)&�D{=��'Y2�w,c	�G�!�^� OR�ɕZ�lSbM¾��tW���8���j�4���h/3}0�Һ&}^�����Aʰz�3L�=:�t��C��r�l_Փ�ũ����O{++�|�-.�d�=��<:��B������E�`�=�����=���%��IG��
�6���<ocf�	"���sɊP��w6W�T%��o��v������>�����"˘/	6�}�Q�����k��Cp��{W����[��oXÖ���b>_���2&����=�b��~(��P �7�r��q�������8���o��H8A����ʐ��-7�|�Y���Q�d�_(��� ���x��d�hKn�
�h uz��y�M��
�O�|7�o9h��K3����&��5��:ܴ�a�6�F�����Eވc��t�D������7�_��-����o����'[N�O�E>7W2ۆ��鱿铀��_�cs~8���E��T��_�(�\К�Rc���S.1��j�V`�"~���e�Lá`��/̸��c���M�d�y�����h��V�T��y��'������w��	�6� �B;�a~-�-�� �zϩ!��b�^��{88���������UϪ��d����#�����H�o���<�O#��K������jvt�����!/��iz�3�젇k"�E 3Zy�dnr�x6nʎy;��$����t��~�9ɰ,`1tO���$0=��@M���:�� �0O7e�D&����h����)������1ږ�B̏��L��z����˾�8�p4�"z[���|��K�t}DpDZ��NN��"���d�ŏ�W���$�w��]�'����3zg�$$eAg����s�Yq�1<,f����>X'�t^FӸ�@�9+á@)�ô4]�^��g��4�l��k��kш��j-�JG��ǐ��P����k�bAKU��V����H�l�W���޲hpmK����7
����`_�h�+d�������/Z.�8"�.���+�����u޽y;�?a���!Ȋپ��?3&���	jd7�	�]�%��w>ޤ������^��op�+M����mޟ���j�`W~:r)��I�*4K;B���B}+n>�@B����I@v޵��o�:{�*q���h�c8�;�O��.�`���.�qxA>YKM˯�췢m:S�:�2���
9~�K��D�0�@uk~M�6�	ҹ_-�!��x7��K�ڕ��s��u���eך�K�b9;VD�W�NcFyl
=��PLlp"��|}y ��2sɈ��O����<�<��c�s�ݕC;*AZj�m�h���Hl��d��34Y|���:^ML%��6�K�@����<1[��u�rZ�|;��GT8�,[���Φ�]E���Z�7�ݳ����xp���o�"������nA���yFZ���g�{���G:��J'{�����"D�����箆�������%��υ�^��H���t�+��ַI����|9�׬�AF������|��H�
�B�IF���~=3��d�Iͻ�������-$����)�;���m:��,���F͝sr�9,\�w��>���	_ĭ�K�G�,弈�<�sm�U*�FL[<3��g��y��]_���_�g&i>�����eL�A�͝���|�G�����ɇ��5��T�����dB��6O���b��T�_@�d��[8��)�	�������[�?� ������Q��!-7R&��ѳ�q�C�x{VR��7��w/z>�-���Ė�m6���`͖����M�Wc� �d�2�g�0������z��E�ʹъ�v��Nx4>��C�*6��Q��� �Ȓ�@p�L����E^�?���z"�#���*}i��uV%����h7lC��4���'�D��^�i[b���0�2�-�}���<��5����	��^r�5 �>$:W�m+䣌��dQF���,��}��Y;�{�e>,b���!��(�/h�����X~�z�wm!��,�يHn1hK�E�-�K]ԃ�Ex��3���>_lq�� E❕�Ƕm��~7U�1���N���n���9m��ٴ�T�N_l��ۘ�����o�R	����?�^�� f�X��o+q�~�ߎ��Ot�
�o�d�p��s���;�T�WB���u/��h����$w��3�ar�������b��6�4��e�:�A����G��ӏ6Ep��v�N"y��D_@Oc�ģe�ytu�Za��xǒl5�C˱oՙ!n`����T0�l���ye�Z��R%�^ʢ<�/���a���17��;5�-�}��+��<�}�>Fֱ?%�J��:�	�6䄮_�<�(��=QNk}�!���j�/��Rr���{G1��\�#����2�V�,G��L`b;�/8��%���X��vJ�} W��4o��9-��5��U����$yU��l'y�������{vL��]7�Y��X���j@_m9�Dp� ��
e/�&���!`i��u���N�!+�㹏x�"��ed�nOo��U���t���:_��oid[�ޙ���̍��z�UN!�J�!��ֵ���m �]�������9刳%�3p2�L