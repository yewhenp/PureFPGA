// videocard_gen.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module videocard_gen (
		output wire [12:0] memory_mem_a,       //       memory.mem_a
		output wire [2:0]  memory_mem_ba,      //             .mem_ba
		output wire        memory_mem_ck,      //             .mem_ck
		output wire        memory_mem_ck_n,    //             .mem_ck_n
		output wire        memory_mem_cke,     //             .mem_cke
		output wire        memory_mem_cs_n,    //             .mem_cs_n
		output wire        memory_mem_ras_n,   //             .mem_ras_n
		output wire        memory_mem_cas_n,   //             .mem_cas_n
		output wire        memory_mem_we_n,    //             .mem_we_n
		output wire        memory_mem_reset_n, //             .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,      //             .mem_dq
		inout  wire        memory_mem_dqs,     //             .mem_dqs
		inout  wire        memory_mem_dqs_n,   //             .mem_dqs_n
		output wire        memory_mem_odt,     //             .mem_odt
		output wire        memory_mem_dm,      //             .mem_dm
		input  wire        memory_oct_rzqin,   //             .oct_rzqin
		input  wire        pll_0_refclk_clk    // pll_0_refclk.clk
	);

	wire         pll_0_outclk0_clk;                                              // pll_0:outclk_0 -> [hps_0:h2f_lw_axi_clk, mm_interconnect_0:pll_0_outclk0_clk, rst_controller_001:clk, videocard_module_0:clk_hps]
	wire         pll_0_outclk1_clk;                                              // pll_0:outclk_1 -> [irq_mapper_002:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, mm_interconnect_0:pll_0_outclk1_clk, rst_controller:clk, videocard_module_0:clk]
	wire         hps_0_h2f_reset_reset;                                          // hps_0:h2f_rst_n -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                  // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                  // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                 // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                  // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                    // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                 // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                 // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                 // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                 // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                  // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                   // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                 // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                 // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                 // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                 // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                 // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                  // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                   // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                 // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_videocard_module_0_avalon_slave_0_readdata;   // videocard_module_0:data_out -> mm_interconnect_0:videocard_module_0_avalon_slave_0_readdata
	wire  [15:0] mm_interconnect_0_videocard_module_0_avalon_slave_0_address;    // mm_interconnect_0:videocard_module_0_avalon_slave_0_address -> videocard_module_0:address
	wire         mm_interconnect_0_videocard_module_0_avalon_slave_0_read;       // mm_interconnect_0:videocard_module_0_avalon_slave_0_read -> videocard_module_0:read
	wire   [3:0] mm_interconnect_0_videocard_module_0_avalon_slave_0_byteenable; // mm_interconnect_0:videocard_module_0_avalon_slave_0_byteenable -> videocard_module_0:byteenable
	wire         mm_interconnect_0_videocard_module_0_avalon_slave_0_write;      // mm_interconnect_0:videocard_module_0_avalon_slave_0_write -> videocard_module_0:write
	wire  [31:0] mm_interconnect_0_videocard_module_0_avalon_slave_0_writedata;  // mm_interconnect_0:videocard_module_0_avalon_slave_0_writedata -> videocard_module_0:data_in
	wire         irq_mapper_receiver0_irq;                                       // videocard_module_0:interrupt_finish -> irq_mapper:receiver0_irq
	wire  [31:0] hps_0_f2h_irq0_irq;                                             // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                             // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         videocard_module_0_interrupt_receiver_irq;                      // irq_mapper_002:sender_irq -> videocard_module_0:interrupt_start
	wire         irq_mapper_002_receiver0_irq;                                   // irq_synchronizer:sender_irq -> irq_mapper_002:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                  // hps_0:h2f_gpio0_irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [irq_mapper_002:reset, irq_synchronizer:sender_reset, mm_interconnect_0:videocard_module_0_reset_sink_reset_bridge_in_reset_reset, videocard_module_0:reset_sink_reset]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	videocard_gen_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_gpio0_irq  (irq_synchronizer_receiver_irq),   // h2f_gpio0_interrupt.irq
		.h2f_gpio1_irq  (),                                // h2f_gpio1_interrupt.irq
		.h2f_gpio2_irq  (),                                // h2f_gpio2_interrupt.irq
		.mem_a          (memory_mem_a),                    //              memory.mem_a
		.mem_ba         (memory_mem_ba),                   //                    .mem_ba
		.mem_ck         (memory_mem_ck),                   //                    .mem_ck
		.mem_ck_n       (memory_mem_ck_n),                 //                    .mem_ck_n
		.mem_cke        (memory_mem_cke),                  //                    .mem_cke
		.mem_cs_n       (memory_mem_cs_n),                 //                    .mem_cs_n
		.mem_ras_n      (memory_mem_ras_n),                //                    .mem_ras_n
		.mem_cas_n      (memory_mem_cas_n),                //                    .mem_cas_n
		.mem_we_n       (memory_mem_we_n),                 //                    .mem_we_n
		.mem_reset_n    (memory_mem_reset_n),              //                    .mem_reset_n
		.mem_dq         (memory_mem_dq),                   //                    .mem_dq
		.mem_dqs        (memory_mem_dqs),                  //                    .mem_dqs
		.mem_dqs_n      (memory_mem_dqs_n),                //                    .mem_dqs_n
		.mem_odt        (memory_mem_odt),                  //                    .mem_odt
		.mem_dm         (memory_mem_dm),                   //                    .mem_dm
		.oct_rzqin      (memory_oct_rzqin),                //                    .oct_rzqin
		.h2f_rst_n      (hps_0_h2f_reset_reset),           //           h2f_reset.reset_n
		.h2f_lw_axi_clk (pll_0_outclk0_clk),               //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (hps_0_h2f_lw_axi_master_awid),    //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (hps_0_h2f_lw_axi_master_awaddr),  //                    .awaddr
		.h2f_lw_AWLEN   (hps_0_h2f_lw_axi_master_awlen),   //                    .awlen
		.h2f_lw_AWSIZE  (hps_0_h2f_lw_axi_master_awsize),  //                    .awsize
		.h2f_lw_AWBURST (hps_0_h2f_lw_axi_master_awburst), //                    .awburst
		.h2f_lw_AWLOCK  (hps_0_h2f_lw_axi_master_awlock),  //                    .awlock
		.h2f_lw_AWCACHE (hps_0_h2f_lw_axi_master_awcache), //                    .awcache
		.h2f_lw_AWPROT  (hps_0_h2f_lw_axi_master_awprot),  //                    .awprot
		.h2f_lw_AWVALID (hps_0_h2f_lw_axi_master_awvalid), //                    .awvalid
		.h2f_lw_AWREADY (hps_0_h2f_lw_axi_master_awready), //                    .awready
		.h2f_lw_WID     (hps_0_h2f_lw_axi_master_wid),     //                    .wid
		.h2f_lw_WDATA   (hps_0_h2f_lw_axi_master_wdata),   //                    .wdata
		.h2f_lw_WSTRB   (hps_0_h2f_lw_axi_master_wstrb),   //                    .wstrb
		.h2f_lw_WLAST   (hps_0_h2f_lw_axi_master_wlast),   //                    .wlast
		.h2f_lw_WVALID  (hps_0_h2f_lw_axi_master_wvalid),  //                    .wvalid
		.h2f_lw_WREADY  (hps_0_h2f_lw_axi_master_wready),  //                    .wready
		.h2f_lw_BID     (hps_0_h2f_lw_axi_master_bid),     //                    .bid
		.h2f_lw_BRESP   (hps_0_h2f_lw_axi_master_bresp),   //                    .bresp
		.h2f_lw_BVALID  (hps_0_h2f_lw_axi_master_bvalid),  //                    .bvalid
		.h2f_lw_BREADY  (hps_0_h2f_lw_axi_master_bready),  //                    .bready
		.h2f_lw_ARID    (hps_0_h2f_lw_axi_master_arid),    //                    .arid
		.h2f_lw_ARADDR  (hps_0_h2f_lw_axi_master_araddr),  //                    .araddr
		.h2f_lw_ARLEN   (hps_0_h2f_lw_axi_master_arlen),   //                    .arlen
		.h2f_lw_ARSIZE  (hps_0_h2f_lw_axi_master_arsize),  //                    .arsize
		.h2f_lw_ARBURST (hps_0_h2f_lw_axi_master_arburst), //                    .arburst
		.h2f_lw_ARLOCK  (hps_0_h2f_lw_axi_master_arlock),  //                    .arlock
		.h2f_lw_ARCACHE (hps_0_h2f_lw_axi_master_arcache), //                    .arcache
		.h2f_lw_ARPROT  (hps_0_h2f_lw_axi_master_arprot),  //                    .arprot
		.h2f_lw_ARVALID (hps_0_h2f_lw_axi_master_arvalid), //                    .arvalid
		.h2f_lw_ARREADY (hps_0_h2f_lw_axi_master_arready), //                    .arready
		.h2f_lw_RID     (hps_0_h2f_lw_axi_master_rid),     //                    .rid
		.h2f_lw_RDATA   (hps_0_h2f_lw_axi_master_rdata),   //                    .rdata
		.h2f_lw_RRESP   (hps_0_h2f_lw_axi_master_rresp),   //                    .rresp
		.h2f_lw_RLAST   (hps_0_h2f_lw_axi_master_rlast),   //                    .rlast
		.h2f_lw_RVALID  (hps_0_h2f_lw_axi_master_rvalid),  //                    .rvalid
		.h2f_lw_RREADY  (hps_0_h2f_lw_axi_master_rready),  //                    .rready
		.f2h_irq_p0     (hps_0_f2h_irq0_irq),              //            f2h_irq0.irq
		.f2h_irq_p1     (hps_0_f2h_irq1_irq)               //            f2h_irq1.irq
	);

	videocard_gen_pll_0 pll_0 (
		.refclk   (pll_0_refclk_clk),       //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),      // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk),      // outclk1.clk
		.locked   ()                        // (terminated)
	);

	videocard_top #(
		.WIDTH (32),
		.BYTES (4)
	) videocard_module_0 (
		.clk              (pll_0_outclk1_clk),                                              //              clock.clk
		.data_in          (mm_interconnect_0_videocard_module_0_avalon_slave_0_writedata),  //     avalon_slave_0.writedata
		.data_out         (mm_interconnect_0_videocard_module_0_avalon_slave_0_readdata),   //                   .readdata
		.address          (mm_interconnect_0_videocard_module_0_avalon_slave_0_address),    //                   .address
		.byteenable       (mm_interconnect_0_videocard_module_0_avalon_slave_0_byteenable), //                   .byteenable
		.write            (mm_interconnect_0_videocard_module_0_avalon_slave_0_write),      //                   .write
		.read             (mm_interconnect_0_videocard_module_0_avalon_slave_0_read),       //                   .read
		.reset_sink_reset (rst_controller_reset_out_reset),                                 //         reset_sink.reset
		.interrupt_start  (videocard_module_0_interrupt_receiver_irq),                      // interrupt_receiver.irq
		.interrupt_finish (irq_mapper_receiver0_irq),                                       //   interrupt_sender.irq
		.clk_hps          (pll_0_outclk0_clk)                                               //          clock_hps.clk
	);

	videocard_gen_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                   //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                 //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                  //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                 //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                 //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                 //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                    //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                  //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                  //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                  //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                 //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                 //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                    //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                  //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                 //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                 //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                   //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                 //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                  //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                 //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                 //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                 //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                    //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                  //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                  //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                  //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                 //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                 //                                                              .rready
		.pll_0_outclk0_clk                                                   (pll_0_outclk0_clk),                                              //                                                 pll_0_outclk0.clk
		.pll_0_outclk1_clk                                                   (pll_0_outclk1_clk),                                              //                                                 pll_0_outclk1.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                             // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.videocard_module_0_reset_sink_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                 //           videocard_module_0_reset_sink_reset_bridge_in_reset.reset
		.videocard_module_0_avalon_slave_0_address                           (mm_interconnect_0_videocard_module_0_avalon_slave_0_address),    //                             videocard_module_0_avalon_slave_0.address
		.videocard_module_0_avalon_slave_0_write                             (mm_interconnect_0_videocard_module_0_avalon_slave_0_write),      //                                                              .write
		.videocard_module_0_avalon_slave_0_read                              (mm_interconnect_0_videocard_module_0_avalon_slave_0_read),       //                                                              .read
		.videocard_module_0_avalon_slave_0_readdata                          (mm_interconnect_0_videocard_module_0_avalon_slave_0_readdata),   //                                                              .readdata
		.videocard_module_0_avalon_slave_0_writedata                         (mm_interconnect_0_videocard_module_0_avalon_slave_0_writedata),  //                                                              .writedata
		.videocard_module_0_avalon_slave_0_byteenable                        (mm_interconnect_0_videocard_module_0_avalon_slave_0_byteenable)  //                                                              .byteenable
	);

	videocard_gen_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	videocard_gen_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	videocard_gen_irq_mapper_002 irq_mapper_002 (
		.clk           (pll_0_outclk1_clk),                         //       clk.clk
		.reset         (rst_controller_reset_out_reset),            // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),              // receiver0.irq
		.sender_irq    (videocard_module_0_interrupt_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_0_outclk1_clk),              //       receiver_clk.clk
		.sender_clk     (pll_0_outclk1_clk),              //         sender_clk.clk
		.receiver_reset (),                               // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_002_receiver0_irq)    //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (pll_0_outclk1_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
