��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ� �t;l-8���[�R����1Bl��v��ʷjϱ3q�`ĳ1��{�?>a�f��,�0&��K注 �%���* �R��D%&�CǪ��ԘH����JK>�+��lM����dd)c�>��N�x񟂾�-U�|9﹉�H8���O`;�^%6^���sb����(�'衄w$)�r!0S�,���y#{s���	��f�$i�YBXZm%�F2��^�����E�Jq�{V�a�����'{����n!&�/���)KM�rN�ڳ ��)�5%O!U���f�:[�� �����mI���a���"�pd[��c�д��f�����	�Ͼ퓮�'@���	o�L/ɱ<v(d��|j(���0t����	��KP��0���1��,K�Ɓ��>Sk�$�����}��g;���c�.���PH��f��O �դ%�|#[�8�-o��n��D���O��T)>�\в#�;���P�U��lN������^�Ҩ.�8��L̴�ݧ�_���8���o���]�z��Q�ӵ��KN�SFl�`|�*��T�U�[���*�����u�XY��	���R�����U{�(����{|���&,k|w�f-��݇��y�޲~���3(Mo�}�����Y��:�?���X����,xm� ���K���)X=Ր-0�:uJ�:~VW�̾�ʽo�3�` �#z��������)�����0T��k��!�Q+?" ���6b�Kn�	R0!�C|$�����j�.�(-���4�,�	��չp��v@�
�2��"r\�de'j媤��3�;p�ޤ�&Uk�e��EU�]�����«Ӿ��@`�,
�`76��-#���Y'"���`��NLy�e�t���D=����q�)��Ɨ���|�ͫe��/�F�?��57As� �?{����x}�Ś��U��c ]Y4��|P_�8�L}���ʇ>�_ ��&�$���?ߙ�g��0$�K�T7u��� �Z~��l[{����Y��R��Ђ!i[�������[>l������ �s��MO"���7���#������y����.C��sy�:���T_8�*���,4Ty��Vo���E\# �'�m>��?�Ϟ��#��5�$Aح�n5��--�Y��R�, s�`�,��E���DgoZ�@w�<��ݜW��Q��.�J:7��{/��.9(}� 
�g��F���vU���j�?\�094�i�Mы����B��
3�{X[��Iz�80. �@��h���N{�z���M��~/��:���wbf�t��
ಉ��[�AVfc�\c�s�|u��z	��Rs�@d�S~M�x�M'Q�)X��ЋwV:��]�k��Wbpq<W%J\T�1v��j�љ����%I����`'�Z\�/�6p�ZwjhU6%cT2����SE �'�h�|V��X@�A��Sf�����6�M��_�UU8g�z�p���.I\�I(SO�o6�=�;�����{�=��NLF.W}/}�@��?
��=7I����e�u��5��k�~n$�q�x������2�W���s^S�C�E=-r��Dm��H䒌L�|@'�Cg���n�[�� ������b�����~ˆ0����՘m��K�Z�E��;�r7US�ff9�m�;���?�]BE
+�6��9*�f�H�t%�2�m�ڼ��sV��#ݵ3���1K���6�TX��^_���/�gQ5���*�L�=��Ա�7�,(�N>zX��[D�bZ����z�ۤk�W1M� �+�_�{\�Mt7/~\�H��<+���x����W�*�ǅ�C���ͯ}�O�f�qW�n�������K2t�pbS�<�c��^��Հ�0~�x�5�w ��A8)%3.��2F=h�I�]�N��1Vy+�'�Q2EɅn*Wв�]�e�Y	j���d�[�i��Y��G՟�b7Mcw�x��F����i֔�1/�����Qf�D������o�1���KX>�������t.*s �1gC��`��$�4G�X���M������X�M�.�s��8�X�6���{3�ؿ�u"�e�]�� �4�_�L�9�s����tSp�;+�j��:�����%{����i5%*�E��������c��G�����=�K���y2���Z}��?�N���G�Z��"x��?�tY��?��FC�JL)N�CƫM�
n
�� MM���X���J�O�[��[2��s���w�c��ZA���S�MGK��c�N����X������g�x���c�!��wɭҜ�ZC�ٗO~icCn�#??lW�S����L��L��O6˙�C5~��rDey�#}LSᩃ�wh�o����� ��L�yC�U&��33�Ϸ�F2�^+�@���P;��.�͙�!���Ǆ�d�I΂h`���pA��[��� /K	� \�X�P!�I��lVk���B�h�u��)(�J���+�kO�����Y$R�4Ҵ!e_�nL������CaW�hd��݂`
�|��L�$��^I"�w�I���'�"�e�w�����i���1�"p`Zd���|�:�Y.��׷b��R���|$�=�G%�Dl� &��釢�{�)�����[K��K��E��v:D��y�ٝ��O2�˓�ҤM���J�wc�~�³_��
�B�=�*�rn5�<����1JA1s����^�n��GazR�AC|��}yOw��t\&+���I ����I><ظ8��JA������r�D���R�fB�4�N�6h=��n���V��Z̰ ���2�W��PO�}ؼz�� @^J)%�M�V���%B@���_-���O{����b���׍�DI���0�Da!�~����|�Ť��on�r�FV��1;�{c�Z�p�@�=Z�)���i���p QτV���$Mp���@&�J�	�75�Q��T@ywylC����,s�]e?�k��(��I�vt��8u9WXy�
̍���aZz�:�M���*�2&�s,��3�a%��c؛��K�>L8*~w{��3���ag��$�������B��S�c���۠�T��n���;P��O2�&R��+��Z�<�Ϙ����\�}����t};�"�����y��緖�}σA;@=]H� aDS"?�C�P�m�lK��Pb��l@�,�a���Ŵx`1�/髣�M9����{���Ez���	���=�R�6-y�d1�~d7���v2����e���B�;f�vK	�$!my��������h4��Z��#��v?;%�y>�v�4��z�܂�f��'���jS��3�S�m^0�!��k��������� p����EG�C?E;|�*tD�@�,w+�V��/l�K��?a�0���ip'>�mc�[�Oz��F��ժ�K����s��!�S�u�	��ٟ��ŕQ�V@��x�A,�w�ٲd,�l���q�fF��@y$\,z�tp��G�#��.o���}V"+�V+��� ����r�4H�Fn�Y#mAZ>��n-��=Ћ-���nU�U��нU9](��T9��\?��Yo��Oy��		*}�7WL�}�Ǔ��뢈r%�g.*P�
	U���^�L6 �ѬA;Y�w-���~:��Ewf�m<����\
���Ї��� �>� T�f���8�T@��w�W����b��h�K�)��OÅV�׊�E����}�I� Cn��##��.�d֝ȍc�y6���}@�����kR$�2⿟yB�i��
�^es�Jw��e��X��U����ĺu�Y��x�|�486��J�K�;����+�7�:��EyN�Rh�wX�[��v7�~�gE��"�X$����w��l"�Ԉ��ME�O��x�vC�פ�,����83u���b+yX�����C��q���$���#c���ܑ\����묳WL�^D 0�%	�\�d�8؂�OЁG�3�%3[kf�e����W���L%��<��F��V$ҡS�����h�N¦�_cx���%Q��x��44�R��?�><ⰶ��1�;(�Ri7�N�ZҷJX#�Ev�w%uevIT���[� ����;�{ِH���&��s�Y��j-+�f�!��S�ä�p����'*�I��y**��-;�-!�S�J	��2��]����U��f�$�}��۹Yt��2�ϱqFt�Z̸$lKA�t���I]������(k��mZ�چ��醻�R�oR��g��J@�Jw6�1cdYU��o{�|N\�6�X�#��I���nm\���{Iٺ��x���%��-� �Nf�Gɒ���{Ĥ����eD�G��+#���a���
R�J;�_�R�*�ħPT+v�IW��� ����C��&�1��L>MJ�&�K���t+V��S�):���,�*Q�"2oMB�����ziU��!�)��!y��J'�K���-��ӫb���ҟA���Ĺ�K)���
øB
ȵ�ά��YhXK�����R�����|�*I~�*s�
�_.���N�wesu�5��Z�:���5�֛�
�C��#�bj�v���'K%����dN��{8l5Q�'#������۳"HK��x���L��8���B���܊�4\�}[M��y�*ss���b�4���cO.m遌�Dڳ��p�"����H�Q�Fi�G��\2��HRo�;�P�F�B����E��l�u����x�P�L������z��/a	i���X�}?�1�Tf�|h�n~N���5Il�j�-�R���R�8�s�V1�����Fs��H��i���VO�%f��P�x��E��x�8P�6�����/�=F=Rd����ٷ�����$�׽a���88ɳ�e���"�S�rT�:���F�q��׎�dӆ��*J*��K�*���eC{1��b�yQ���(X�^-/Jm�W5\��<%�����g��KN�N���eׂ%[a]Sd
c3a���B�7�Ff�N�"��
:f�wE�Z9����&�b����{� ���K�q�p,��l��� qMY��:���
�`�L@55mr=�J}Bz仈�����Z
�@��(8P��������H��6�O�F�T���E@
Y�n]e��Y��Q��t���W�ү�yx����Vbحڮ�?L@s��|���O�"��U5��X����ׯ�/�NN ރ��Vf�����Pܳ�w	94�24U"��P�0zm3%�E�  h���R����W���AQC
�+m
��8<�\L�T�yW�G�4k�"�ۖ���}䏑 �;ӑ�ߺ�lia�����ot?`�&�;�zi@/��]��`�A/tF!�_̍������T��lR�ډ�&]mނ|�ne������4oG���M����~����|k�Og�^���GKD%w_�zn�C�i8�ɏF�A�#���M��y~bb�����23�r�zDr'�y�U���k���S��H��CC�D�М��Kɉ �"צ%�~qm�#ڲ��X��7��>lߜ�?�|$�2�ނ.�.\��rU�$|�K5����K2�����_���n�'��r�n�ė償M��>��_|��*����P ��ff�F3l�&
}!�O\�+o	MR�J�c�l�<���[͎�8�kܴI%_nHl��7s@ơ�@�]�*aC�\�T�����^�`��|�8�Gʣw���3����Ӑ-�R���e�K��xA	!`J�(@�0B-��-$���p~W��#�.�t�R��1�|C$�x
a�iPF���h;́��Z��"��ޚǨGʬ���S���H�'��?��)��8�;�qt�Z�@��R�H4*D���;~���,Y0�f+�Ac ��`�u�Ռj0}k�n~�R�K�sKg��j8���R?� ��?�
J�%�ԕA:�&��Y�v���g8�9�������p*�{X�+���e3w2��B�i co���}ub4`=�}��䒿�$䃋�q�׌-�f�R�]�
_H�l��u������Qϓ�.�ge�N����B�~��n~&�i�nY� U�N�����؃Mv#��b$
��l%�.��KzQֈ
�{��5�d�*� m��M�YX¯*�x��-�X)��n1}�����ԣ@����l��!��x��5(��^[B�[�Wi�`[i��ə���]�撅�Km�쫪^�[�7�g�b�ׅ�<hR݂��Y�|��	0)?-�N�������LU�����9O�1��<5�T)7�-��|�}��T�v����Ң�@�+;=x�7:�,#��1�xcCA��m�Լ�9�"vYF��J��ے�@c0K�WBaֈG12���|���X,��m�ߤ�㝩�ۭԑ���
�� f`�����~�3�i��<o<'��EN��*��GV$P�=��ځ���7���pPz�Q����L��əE��j�hќ���f�rN�ó�[S�(h��U�Iy��SY�=�0�&�z���)ە�2�Y��O?crq�	���!��6��4<�o�$F���!�|�{L�e��@aQ�t�\
���h�?~(̳
���8c�6�����GfQw��lbx��Q��%�	����7n�(��PΊ�(iQ�?��g�ߺ�փ���>S،8no=���y�ӣC�LT�;'�K4�� �#�3����0����Ma��]��y
���ЉO�C&� K�n����~�})�)�!w��^�a���r렊�9u��tg�;C�GX�L���jՖ��H� �d/8x��~�I��j9N����xA��T���{P}�ƞ��:��RS��Y�u���͑Cq�D����~:���T"�%�l���蜏�&:����|V�54���:�ߠl��d.��`Dn�"�����]B:�wjӃ�|W)��f��6��J�Sﰖ�fuN�UAǾ{�6v͡��#��2���L/�51,�@��ڲ���n��lU��|<� Q�XW!?/�a{k�|���β�:�SU`ywz�<_�?,Mxe�/�\�C=!�%��:o��q�,�.;߸G�ɋB��Tϰ
Q<7}=��#�oޜ�+2�G3[A ��5���'hEYM��C^�IDZ~
(��KU[�y2}�9�0C~��d��\0��Z5�g-	ی�x�ū��\M� BrHv�
Lm,�	�Hi%���e��D}\��� �wzE��˼0z\�&!*UB:���r�w�A�#����H�,g�3�
��;�<'/�y(l�n��������l8S?���>�S��07��B��'e��՝�p���� ��&/�Դ������J�c�z��<ͬ�c�H+�$1��t��͒i�����:�܄��(L}��i@�*��401����T��!E�%*���P@A��P.�Р0*�F�/:����=[r����o,�"��"��\�7~aHM�r(F4����J�& �,��+��6��:�}cH�0�N�pL��K3����J�
a�a�#� �gv:7������i��(ǝ?+O5�g&���?�x�.{,EnBB�~8TF�v��
�@��g�L���A�;{�<bu_:�����G?�D�5p��W�YX6�ώ�v��_'�q	q�Ѹ�2�ٝ;hQ�&{�K��&����W�}oiٗн1[k���ʐ����{
̾
o�A�.�%\�5�d�E%�a87��2�ּ7ݩ��Rh}���n���0,dhD�}���.���d�s�Lq�Fj�y������:::UL��I�{��g��6��;�������SC�XZ�?�����a!��Y�d-yuܿ3�C�D��	A�ETK�ἄ��l��[a�?.LKI�����hheb��Z�$�y�K�}~�,�j���Z]$Ån)p'^�3X�p�Ù�ut�M�G`�*�x3��i;�S�+���4x�����z�1�{�rH�T%�J{ш�~���팣�8z�Ie�V��}������ս�����`����zԚ��9T46��)nځL��oM3=:# `���m����"���� m��U����k@�mJ��3#T>�$V���@�HԂ1��S�e�j��� ՠp���oam��R<�O�Ƿ�Hq@�8�s�[RW�@�^��M�%�gJ���i"������bu#��?��yѬ��>	�l�Z���y�u'HTL��'c�cc֫�R>�!I�I�ݗ��#��ͦ0�2=9z�#Ͷ#���*���\�Q\m6�c��Z��Nvk}R��r��9�t�Fe�L���}3�Ys|*�y^-��� ��!�`��ۿ-:=���/A�h�a�͓��=�� �|1��;¾�xd�"� јh!$"��@LE�ԍm���F��Ro�ƭ�d����彥v���DF�g<��i6f��dæ�[����`���ҍM@<M�9|�����l
�]U(�֢�нXx� PbNw
��E�2]�[d<�wR�� �i����\7ٽ��{�o=�\Ɖ0��|����K�R��f�k?��Pz��]�1�A��j�/y�O2�\ ���2�#,�H� &�B��}F�7^���A@>%kd����"(�!1�-:42��c� ������#���qT���������`J��q�$8v>�8Hb䤘�%��5�8��Q�0�7�HeT��<��7HXL����U~���
!�Y���8E8m��=�u���R2k/���mۏ�%YTֺ��zB�/�1��gח+<}M�~��ȧ��z�]���+Q���t�xo�qƴ#��n�S�a�Vަ=5�$Ў��x0(Ӗq*k���M�Q�����k�::����!g���+q��7:�Ē�i�!��,�6j �]C���?��?��i�e�e��s�sӖ �@ 0����P�٪wY�q.�%Ђ��
��eQMs����c����4z'ELq��t��򩢐%�`�ιp�q��TgRe����#�Q�>[m���7# ��np
~CBB�cǱ����y���:yy�(z�b0�ƨ�8�	��Lk*KB	��)�~IE��6qn�YT�Y�S��h0���{�	�q��E ��>(IWY�D*���c*����$�1�Mn���8��P\lf�S?�����y7�1\��f�P�X���P�z��*9�4R �4lCQ�oGl����f*xM�� �g�D�r5�������h�	�0/+4�U@u�1z�����ͦ8���l(Cn~��e��GG�ʵ=?x���ɇ˶�Nyh�J��:6_�L��uX���o�JT�-h`��äD��A����Z����s|r�eE��cG�Z��E]��9��0���i���d�F�HׅƳȟ4��gq�V�q�:����WMB%+����'���*s��۷<��Y�Y|6%7�O����;49�)�Ş@#-����>�$�x�ȁ���zF��P$������@���ړ����X���j��2�,4���'�Ѱ'���$ʌM�jן3��M,��<�z�Q�|^����b)$���af����TI��{ ��se��ȼ�e�o��M��^�^��E]+l~��&�+�vCX{�{�iF<��
���H'>���F�K�d��)y�&A���a cn`Ob~��>�F&��$��U�$�)!�7�\�xqPWc@�"�*~��i�n ��{�',bҟ
U(-��3X����X|UV��9����I{!�x�D�A|ֶI�O��Tff�Pܩ�N���~#;w^y
��$:2�W|P�h�@bFtA���j>���Y��mdW��q�?�����*>� �`��*b��.]?�r���[�ɰe��-�JӮ��|�������7a�讴2K�����Pl���)"s���c��P���$��M1���]�%⻰z�ڪ@��M�2Q�I�'1����C��|/m֛�v���*��q��M�rd%�־�A_���"�!�^=-[�.ܾ7�dɣ�=\�C+�����EД.Si�Omj,�g���3V%�4H�"��wXr��P�Д<eg[:��� ���MG��=�Q��%��D�*�g�J�/K�c�ZL�t�MlԠx��{r��z>�MR30��'f�Yr�>,�^I�5���ˠ��HcK���	��N�V���x�",P�����Ct����W3���K̋�I41�E#�(��)Eo���:DM�M�N+���������ܦP͡Pƶ�?}��4�\�W�Jܼ��R($��1EL`�d�Vߔb�M��ܤ�[��/�Xʏ-G ��
M�ϹL=,���-0��?�X��W�E�p�wp�NgD�b�l�e�^�B�q&�B�"�*��*S����I�x�"b9<��@\;��!� ��JFe�D�e�W%�����:wV�vt�q�p��'(q(�P3���7�.��A/mi��]����M'�d��/+|1����4HB0���)����3�F	���u-�u�*������9��Ǽψ-E�s|��W��$�mkq�]�lM	+��`>�Kb�P��q@�`V!��ꛝ {�MIE/VC�h9� ��%�#�ޘ����e���J4�L��9�vq�ߣO��3��G|�vJ���\�94�H+Ѯ�5�?~�����
�&��,���P.�tɲ��xX�
�J��d��6P.f��vN�:&19�A��~��åd���O����b�W�<Nf:�n���i��y����,rǲo\� ������>bO@̟�D��wk���q^%�,ò���1#�Df�����9`��ʀt��jPǶ�`�H\�(����� $H
� �/�D�-���=�ScR� ~�����:��/p81T���D[�0Ļ�g�^_~������.O�%2g�&ۏ���Z��^���9ce��;�z��ձ�=����MG�|�T2L� 4��s����]?\>�����gט�l �?j����Uq�V:;g�ݤsye�cC@Z��L��7���x�N��2�p��78~.�ɒ7V#��Ӆ�z.��WY9X�g*�Q`��3˩g�FJ�I��4��0�
��ֳ�l�cN���@�yz�Lԥߖ$���u�J�-/�^U��v��Q�\<�1�=ao�%P�8#����}P��"A:Z�q�o9 �>+��]�)vM�І�[i�o{ܓ�1;�O�@������֎S��XZl�H�6SU�ۺ��w�VR���-+;��Ef��d�?��`�V=R��I�h��K��;��-(��yy�����x��ES�ᡫ�����%����I�.����N��~=.Bz����fl]-O;P'-M��!Fc�-���.���E��%�i7�����9�
�Y��dy�a2��#'7��)�� ]��K�}a�Ҫʪ^�l�uG�d*�j)%���(8�<��}����:�+�ٖj�.a��p	%o;0yգ����U�RM�k��$�rņ��m)��MvA{���P���e�Qg&���w�N� ��l�abDk��4�!DX�`��2���7�#8�,�]W�
`����:zcm�X0{9�Sc��&�S؉�0y����^lbŖ1���|�M���U6�iW�A���h=�%�0�-E)��tל���;�X�����L���
�P|9���xg&M�	���^=]#e.�x4�yg?|}jaͨ���e��.�{0<�~6q�B���\���x}���4:��	��p���$A�'�d`U���hN�`�}������8�w�3�
�kk\�1��vZ�!��h4#Z�\�t�~��UZ��ťX�q4���rI;�R^7N���:��MV���!+/m��{߹p��W��6�'qϒ����#�La-ʉ}���~9MQ/�4��x�o�>|5��"*��m �?���}p����#��ӊH�c�mȍ�sG�p$����d�m�U����;�jB����>%Gu�_��d9���y���(/��$�b�do�x�7����`��p@r_�8,�d�w�����=9�.�S�� T؏l -�ȕ��2�ߖ�##�Y��F	�5ls�i���X=cA��T߄������F)�wp�mS���{4qP�[���$�ak,�-�`�)uyb��.\�ܓj8���_���ݨ�����VR��$G����� 
rt����*�2^�s�����Z%I���v7�d%�C�>lR�B�t���J�$겸U��(u䨑��rkuH��d��[<[��y�{w�J�p�-ɞ�aspޠ�T�LD�0�@�r�D3ׄ�ev�í�~�|va*&+6�b��O~N�����>{�� )"�4�q-���3$4H���ۙÀ�\�{�'�&ټ|�(ض��пf���8<��M���3��t�~=_�>��{�u�4�XG��)m�.��4$���0F��e)׍�-w˖^[�)
���]:���?tw�}�/P`:ՉQZ0��W���Fe	$��zB3��=|�ixA��P>�|����Gґ򟢾��4�Ř����t3_�,��28~R\���-�]������Hy��N;Tn��6�����5�h8=��'��Q������P�v�
[W)k}1;i;em�8��,�����|�;l�L�X���[�����ѸCL�E��f��6�~�I���	Q����EB��UV��1'���]��8i�v�Z���8���k'�R�Ӎ
����*�JR�8쵃_s{���~社S����Y7kk]�0t�$�ʣ�&O��I��=��5a�7������Ek)O=6�>�!�"����Wi�gI��Rd6[��u�L"��'���;�QU,ryY��:��'�����]�xR�����"Ll;gd8�q�Sla����S`|�m0S�Ǣ�p������U�~�0aa�����y�4a69P9�Sba��BI���"��I��Nj�T`2�eW�U!��0�aC�����ޝٮ�W������J֥��yFٱo���{}|R�[ K�C��WI0�9���,��6�Dj�7��t�A�ac������Z���\�SR�4�2̯�^����ԛR���ȑq)A*m���p.W��������B0�혀�@��<�r4���t	��-�W����  :-��hl_�%��� ���X�v���m���0���-����6�
���p?�A��Bp��N|=-���y����1YE9�![��B<��P�����X�/Aw�Q���%]��j��c��V֜5$�B��?�Ɉd�㶠>V h?e�3�,f��H�l�U�`�n�m����q���1_��V��)-#:c�H�VP�g�Ξ��L�w�&����4p�S��t�"��Q��ϸ�����bE-jQ�۾ 3��ܶ�Ԓ��� #<1��~Ɣ���xzo�x������E~5��Wy5�|l7�E�&�Za� �\q��D�ہs^$�S�k
um���C]��%I��P���o�š�h��U8�K��ɿ����$1vY���a ��M����$\�l7�DF�etR�012���7h��Js�%e���|�Ǉ�=�o?E�"Fgg|� !!�'�~�gV��!M�"��6��*� 3m������1x ���-[I��b��(�!��9�'�8�C�hhܷ��?&�r�m��6ۉh�8�#c/�o9X�L���kjց�>��J� ���T�� �S�6�qd����c
��X�(�&� �-�����!*���Ǽm�i3��m��pOwc�ɋE��ʞ�j���`L�曌�;�Phїլ��\�AM�@�(�;�~�v���ӵ�4��F�#bq+�$��^�*u�r_�M}��*F���t����5����X��^�n#�^x}���x
e6Q!�z{ds����?	��l�ߋ0��[���� <.+�F�;P3_�c_\���Tz\����.�Y"Y�R`FL�;��9�U�(�=���j\	�ɟ\�`�܌+~Iu�'���+5�=���(N�~��,,R�-`��j��>'���S�P�7����[��Y���?rո���.���Q�elltY~�+�Z�-/@��8���������z����}�P��$�q���";"wё`�dS:~��\��O��c���JΜ.��fls<�o�GԇK����̝�@9C�����;��i[�_���@!�~��q����4�5�T>@
�#\�6?���zi(�����%!��[�̾�߄�Z_�;�6���u����.f[��`��k���*�К�d�!+/�I�fT�AejR*��*��=B�42hێ���@�{�-�	����G��('7[�#����&\gQ`�-]pϘ����� �ɣ��UY%����o���45���Ť~��\��%$� ���e`��N�&?]h$mB@8�be�8�/^�xi��08'��Cpf�d��t��/1`��[�:����в�Wj����+Ҧ����`����\����*�`Z$B|V^ujgr	_+<��1�_�~"` F�Åה"��P� (��jA�߶" 7����=:
#���גV�w��m'�"�!V��_��&ʭ�U�N�4�M�鎇�l69Gd��4u�,�N|�]V���&�)%�9�DF�=F�e()��L�����U�$����vv�0�GU��l{�Vc��7���6_��iD���㙮�Ƨdw���T]*)�a{;��+/��0	��:ژ>�^�(폎������6�{�@��A=��9Y���K}/�el����C|u����� I�UMvTy�N1��7K<LE�T9:͗�(zC��3�C3�ˡڤ���0ej�_6w���[���^��k ~z�oi-]�a�|3��<k����1����k#���Z�<��J\�����]��W�D�uU
	�;��A�.�����Q����&�!�OW��W���y�N����b�	�U��Y�h}�˛��e&G�u����<xg*���_�`�Ѳ����F��j꼈 J���Z>f�Z�w�~\���i����
��� ����H0������� �wl�TΠ��0�j }N��<F2oHee���?�4��?�ʆ֘�gC��&���n!���D1�d5��%�nX��L��I+��B��z�\[-	�r�����G?�@�OA�fz9a�V���b3i⠔^*_X�Ub�t��lUz���z���K:[3����D��K��F%	���]m���s	���
)��ؠ�ĕL��������桿]�)2~��VE������썪5_X���(����L�C���*�O�	8v1V����6o�[1 ����?S*��Tˋ�����	�W���C~�2�Yr!�M��$A[6�O��bq��"oW�������$|y`���\S@��UT��)�Y�*�f{����A�CD�;E� [�_�b��l1��j�e�#݄Fv�X�+@	X[�>_^*�8#:a��:
)�,X���)y�Έ��	A�=3��R�X<�j������*�Cy�hjR��[�}?��)j��_�p����")
1�r6:�%g�Ġ��!i&�Y�{�Jv^�f�~-�&�ld���f��c-F����J�&fyl����픇/qk�;�
I�P?I�S�f)C�v�m������珋Gzb�����fH}�|N	Iնnc��s�� 0��xڛG)��I�a.ٸ~�m�`�s��\�����g�R�s�D��L&�E�O�M���(.ÊxBHL����%Վ	�?Ʈ�nA��j�@|�<���VZK际��n��..i�#�C�d�����v��e���hOm�����Ɲ�F .P(��58�fu�U�UztV���T4N������q���
Q&�n)8=�F�~t��v�a��d�F3]�F�s���k,Q�>-��|�:���>k�}��cV$������C�@s�
����J���گ�+�lՏ�0�%��,��p�T7�D��5RJ5�b�j)�V�h�L�F�S���$*����Z�	������X��k�Į��N1| �ɣt��,�WrKO��,AUí�����psT,/̍3�5���Y6�Z����S���'�-��ӫU�Q���8$q=r�U����g�mx|z�w��x�T2$K�"�lZA_�O�`4�,��XϿ�=�ğ�<���4;d�/;��ݽ�sg�j�~�P�[�B��N�@�|�P����⹑���9k��uOFQ��QhI��Uo�Uy����� .3��ҷt�b؀��e̠�FE6��>`w�]��*mO�-��
���j��Z1��<�ç�% V�A�P`ly����ᴧ�.��	�f�3��*��0���ҤuD�ju�G*.pc\Qu{�p�*��tR@�JC"�t�_�)��[[.ٱ�L�����G�������{Ú��)�k���m��H�B��В�/V�X~�=��6c�̝�Ց=4s��}�CT�xuA�w2I����3��:4�y�C�?��vS놋����̄"�|�h���"m���%�@�D���$PI�f�1�� ��gП:2]������Ts���*;}N�u�Q�Xr�NtВ�s��f��a�|u�0<�#��2ŝT�ݤ��EE��A�$tzA��n/M��V�+��a��w��N���zlӇ���E I���j��9�p��_'�fq�'8u�*�����3m�6�S=��{Kb�خ�]�^͙m�������;��+x�yW9��Պ��V朩@��h����vr�i�i��D}f��6����a"��^�q;�m����wL��=�)X-!���a.�3�E��GQ�
HzQ��%��$�s���a�_dîR~=�\^�}nޓ4��e-Y�,�Rx�b��.j�55Z�X��Vw�.9en�A%D��TZϝ~�`[Z�i)�4�!gǐ�kma
�]ǵq|iv�f������W��&&�r�ף���I�<s8��&��A&Iy�e��}ײ�gE�BZ���M��KC�����1k~���v�̗i��g��X�E����=ꈅ$�OY�޺��'�)
&~5,V���V(4�2����f�u��E4����4r�Y,)1�wK��#��o��1{!�ܙ� �X��	Q�
)���ܕ��RI����O�>�v�%�bJKbՎB�ڍ�����0�	s�[���8�`���_=�hw:{�*f>������0-���� �I��6i�\�y��J/1�f͒}�����ҳDѯ.�A�$�{jB$�EM���C	,�����ђ�5�� ���ȥ�0�"VvM�>�L�b�'{/C�FW�e3��>��D1F<> >yۚDg�ǖf�+��Ә�ċO��j��⡜<�G{��}�z:X�$5�ƒgh��ai����5^�'��k��)qԮ���]2p���yR"V�����OfN�wc:ZX�ˤ�UA8'�eΤ�����1�W��=�oNupp�Pފȃ?ж���O�#��cPl$�-/�u�Pz�֙��~�S��^��(��`�#�3E���;!PeLd�#�s�D�~=Xї�Lk&�s��3m_ڴ�^u�3:n�"� �i�.�k���iTׁ��>S�F�5��YMS9�n'"?8؄�qKȫ�V.��β�P~������A*mzLU�݊���z|z0�e� L�6+Z�������'	T��4 7��f17	���&�|̩�P�2_�ʽ��L�,:rK�"3�ȭ��z��r����;'{5��LY�}�(�9*:��z��J����گnѠ�6��Ʋ�Gl?�6%Δj:Eǯ�<�1�;Vc�Y+sc�z)x�8�ا#�ho�yԞ�p���_m�}uZ��;	��`���_�����U�R���b�ʦ+��fp�;z�V��9��퓷��s&�vu��,9P��Tː��H� ���RA� ��O�}�RY��)E�F���<~3�y�e�bI=�"d�DpD��B �ib��� [C��]n��vf��I��Fh����i4����+k��%a,��'H��o�g�fU�!�ԉC�WZ��������̃�?n�Y+���z������v��Cmu�rM  ���q������|%4�7zNDo�H��J9��$.��jy{Z��tʝ�[2>�&����E�t����Cr-D����sn�Ǉ帄O1�f��BE��N�>����5PK��P]��o���u��]�g�uP{���x`�"ˌb�h��P<۱9
I;���N��75�[ ��8Ԭ�ۇ.r�!�{�[��2�J�K���S�`�G���$ݰ<���aóu�;A�%���H�;/�(L}�F��=6
�W3��C�����#�[��Y��_�`A�G��G�;Y����@+�'��_�v�N(��!�%��hɯF:7����"�Y�_Q�CD>�V8���[3�U\K���u:�L���̮�cO�\���f#��݈��y�6��‚����ʴ�X!$��]�aaO���x�6 q�dS()2["�����5Gn ����� y	��?�I�0O �&���:�iS.����}�[Y�����������iOHN��3�:h�>zn�-*3���E]�K�~~�1މ)}U>dԮs^T���Mɺ��꺹�|�'ea�m�q��
������B���<���i��5!$�P�B74.�!q�b�Q ֐�k�ȝI�z��JHW덣E�- �1��ʒ��b�G��d�C��ș�H���"��ŧ��]-GcH'�@T�qo �T������ĉ�
�_GG ������j&x����L�r�gϓޢ�f�C�S�ь�!�,�hإ)%�A��k5�`��<G�J���3�,�M*
�0�z�aI9G1X&:��[J5x0+�D4��ȹ�.�@�-=��p��D휯jZ�����J�T�eM:B�}Xk��ii��Tn�aQFiP���,�`z�enf�v�G~��
��;�<�,���	�㍻�8K!W�F̒/�VȎa�x��1���4K�Bl�pd��+��3�c����GW��IpA�X#i]y6c��t�"aD����"2��4փ�I0X��Y�"\�նb&+$o�5��)��������4o9~/�!�d�o�=Wj�dx�>|��uWK�MZF�s~�
��ϟ��WD�П��3��jߵ��,�����꓂��lV�c�t�l!Vf�T� #�*�E��2�I�=�/\�8o�U�s����+YRi6_��QmN�����>-�l�C)B�zd&6b���Aw�ď�16�M�d�f�J���3N�,\f	�M���_v�a^KW|�����s�[mZ��A,�'�>�����D���ZN�5��ݧ)���ň%���ȓ܀
�9��Z�lFJ���P��|~��,�7��n�d[�%\R�4cݦ�=���u��)�u�G�Ǎ.�&��>�ݥ����3���`&�cb�a��R40��l ����ԟy�Ij I80#����{�Jo�Ou/?�����dG]/=�C�᧓$�U���*�����x<x�h"����(�j �kp��q�9�X����0I�3���cW��c�m7�x�ϡ���+42Af�霺T�^���Lx
[�"�_�����y��H�І�(�D� Mi␆��8<V���"�uÎ�'�[��e�ITK��C������]K@ݓd�|�5�9z�H]��nb�w�?s��ӹ�KSasJ����W��W!UX�'�)��0W�i�xn�{�J�!؊US��o��Q�%��+�Z�zK<T�:C-��d�3baU�Q:eq=����s'�oeI�s�η�������k ��:aS�n����yu�C(M5V�[Jx7�A=L�$^2��7��؜vB=U-��H�u�Y���k8��+!��vl��9}^���ʷ��Ϫ���6<����ww�t�[р��N����-��"��鴹E�(TviI�̓�3�U���(�t�O_3����-�5E�Ǜ�0|m�A�I���٬E��>�@|"�6��Ư0;1�/!DPx��k��m�,R�+��h�>|���īR�_^f�$/h���E����a��}��<�Y���`�|��Ua�����E�t4v��jo 
�WF�C�@�����o�v ׎����VZ*a���d�U|��}7_���o�i�IU���X ����A�Ph�o���դ՝��A`i�
<غ�����sM|��ek�-�-A�4�x��i0��f�y釗���:����|B~�% �`���t��8G�ht3�O�W���D��	{wO�n%Q	y��76*>��㜄in�K�:��_$��h���Dd�)yw����9�o�.!
�oNPAuvz��
����C�O����3P{����/dr,�A ���Z�}�nh���do� ԩP����sd7���̥�<�����)O]tU#�v*�跒z?d����z�XL�v��N}�1Qt�՟-1��@/Z���8��m��J�F��XD4���J~o�7����e-�1ٚ���ʁ̯�%c��a��7Da���q���EE	�_w�Rp��'�RSϟ�D��(�>�R�w��uj�_�܊����mݩ�b��E
�`��T����-�ufX!��n9�[�7yS�����b��A�H7���*��� ����B�ѳ܋π=�cTK������:U���c
��o`���L�s����.~��e���KV�>K2x���UVJ�w~�n�CG���`�xu��ю��v����7���w����k�8;ש�/`���0��Mle}pf��m��q2�$O4ONY�dϷ���	��	%�ׇF븍�� ����ta.w#z"�i�-x�*h�B޷�[^~9ҬނI �T������2m�\J,�;�u�a�@�֪��$ήHK�Y�@�]�W�i��n��&5�!mW }Ms��,=��g���;�e�d�p�v
Hy��̎�}��� m����儋�/F����5���X3�Tc��,�~b������ \Xv�`���&]�m/�5��𿆹��?#?�m��ע��6-��Y2B��#*� 6
u�r�J��E�iXN�[��̧�cQ�\�M`ktݾ��^��"=n��L��4� ����<n��o6T\U�<�k�x�ǲr��]�]��sV���ʙ��l'�k��Q�����d@~$�~�67AM�M�3�M��`��|f�!�����rI/h��4K~���О��zQ�N�2ih��I�����{wh}���WP?�v2�tq�YgM��oj6�o=��0͎>�d�~�ƕ,�}���%?	}%խ8�漵5@k�8���}m��vaӅvU�C�͝���1�hs����&��ٰ��|"�*�>:����ӑ�uݎ-yW�`U2��R�=
#��Ȧ��<��>�O�|'�=ة�!����9ꝍ���>�=U:+>iƂ:��6aD룴�A��g
����w,Ŕ������(�c� /7��铨�Pɥ*���|_��6u���,�3i2��0�����iھ}e�;V.�V�Nє�lD����y��9^�����y�Ⓟ�sJ�q��,�x��8�z���r(L��\6�ժE�
����O�˳�g����x�&�D=8p$��VR�F����M���c��}='M�� ��n��߳o ��$ɛR+�g�Ė�@,���'pe	$dQ9�N�)ҭ=��ͽeC;��F
Q��1��`��rc�G���-R�/>�e�J��2����^��9��
�7�Rߦ�!#eb�&�*K���" �2f}�6�o�D���ԁ�3�a>q��<��(g�!k7`��2NRomP�ԗ����]��\�Ra�h���� ��T�u�=�IG
���q@4���PF��+C�Eځ��ks��Gt�'�c��b���gg��V�w�U�y�����(���W��C6�c�L�չ]u������`]q�m�9��L��[�	�CNdᝲ���V��w����S��6n4&��9f
��iC*��v�JZ�6����^���xKi�o�;�����3�!#��	y*v��~���KH�?	�P2��!O�����CGz���B��Z��%��H0xW� 4�6Z%k�B%uף6U�JO����oDLDȽ����{�7���ܔY���z�a@r��k��6��3�,��vY��6.��Й���^��1Ɍ�$�	�3� �S��'T�����[�a�Oiۋ9n�f9��0�{��5�c\�K��Ȫh���` 0i���>�Ҡ�W��z�X5��5�xB����;0c��/�)#��H���7[�� 	�൴�;T�0 �H��['|��5�$��kW!��K]
�G�o]s�a��Uľ+�O��yT�i���mkx:�j���+�X�cG�+��u5�N�K����`�jA�tf�y��PK�+[mW��N��]R���f�%�x�=%(#1��'�hT�$�@�|��r�iX�|�2w[�,�z6LV.�V���'��̌?b�َK㞚/!�G���f����6�rP��"���чj$�<��R܃��JQ���@)��x�^e��k+W%:t���Ʀ�N4�Z $�?O�����[$aG ~u�-�=?�I_]^P���83Hre�:�h�89S�
4��R�nd��zEh����M���Qc�,d�[!�y��C�6O�i� �;<��$V6����׋�.�g����c���~�$hi�*u��W���d-�s��=�p2)�Us�Őm��2Zyra	7����Ƚ����ʞ�=�~�G�f���#��%�R��	�U3��)]����Xݦ�Õ�m5^�f���uJn�c?�n	,�Z��خVh>գV�����(�xIl��>/R��R��6�@N��y�k��D��>����k8M'��,d��Mu����y��XUq�8��lc����p#���uc����������ڛ�=��Z��(���yGyf���$J֕�w�:0��u.�@����SID�`�S�� 3ֱ��6���7�#j�%�O�=7��9&�;�8�Wq�=���Ç
����������}��&�S3������3�������B�$tB+�[*e���0캱4Kq���5�'A��M��@ Z��pK�#���_���b���=����D���7Sq���+�SO�Ԁ~�9}�,��[Rʧ����xY5�xJ��?� ���b�	� }m�C��Ĥ��,�D?ϸ3՚M<=�pWU�?Kw�Ҥ�S���\��#ɍ��(�r��4��r��7�6���� 3��{☍H
�o�1㮾�T>�z����S��{p��޾����vҧ�U���Z�h�"&jc�V��1��^h�u�g�9�i��N����5W�?�{��a�t�����Xѳ�9�|s	[��42��#	B]Xp��Yp�5o{Uu��ç5t�N�S�o���"����E�᷅u?cfv�;���i�w�;^,��g5 Q����|���h������^=�cx��s�p��A��w=���aX���b�Ya��G0͡ve`�s�Zj�	14��=#s�v�9t=�;���v�Ir�T��vɒ�%��}�::��:���<�(ҍ��R����o�b�VT01�)�̻� p;���p�qU�{�ڥ�o����ڋ�v��aB�% ���"��+�4ۣ��������o�����j�I>;����.�61��n]�e ԌU���T0��3���R�Gu�!�U�W�� ��2`9lׂ��%U�Յ����g���Η��g����8q��U������H�4��r7
��|�̡H�����3e�j��#e���]xHr�wl���h1�\6��$��E�����F����W��(�hі`��W��=�F�w�m�"7x��= ��٦��G���\s�k�"h7ui�՜O�LyD�ss�J�M7��ݴ�F���P�`%�����S��7�Ԑ@�j[<�s�������g��DFD2
��/�B�t�x��#�WV�R�{��;QU8��s=�>��̢������ymۉ��w�;.[���<k�i)��)v��3Ǘ�^D�:E����k
�H�رٲ��M;|G�Ѥ�A�Ϧf�\��կ���(�v�v�XQ?�=�b����3+���*��u�E���~ץ6�H�]�3���aZ=�;py����#^'9ep��o�?��(M�9����=�\G���������_mRa�Fy��9��Ҷx��؇�u4FScN2ۈ_�Kg���W��%��8WL��%\�R��|�7����dR)����#n�x�E<��jc�L9��nN�Qp:Z�Ug��*X�y�ao��=Fi��M��,|��-"�Zi�\b�,��"Hi"�4�a6N�Qc�C�.��Fg]`�x�<���SJ��m�V� [^s"��}�����_��x���[�k�$���K�L�Nc8��(����>����g�ǬP�y�7\�����vE �򚚚i*��r"L�x�� �':k���H���ֱ&��A��&D�T�myH�?�n�M���'"M1H�{�O�'��`�3���7��>�E�Jb��� չ��q�}�M�}���$��c�O"~��Y�{f��w啖��a�Wr?���-j��C]�AOE�m�@H�Qce�X
+H��vݯ�D����i(��㽶�a�M�$_��9��w�����B�ۛ���鸯�VX�@�f�x�@r�W�G�#~��jaA����'y��;����R��^�$�ެ�?�{��8W;���\׸��?���n��Fp��(����l/�9��'[yuSY4Q*��piS����k|�[d#)| ���־�����T��,�8���㩚�t��m�Ơ���Ȇ��#Ő8(��\�֌l�fc����G4b�p�4�IP8�Z#	�մo��ĩ�~�^�ˠ)��Pz�w�1�wO���Nd^A'�#�iDݺA�k��I�",ij@ߞ���~=G�d�5,*mpfpj4dD�v?̑��rX,���J��/X�f/��+�J�t<C��v�5��.�5�ݦ(�1������à�H�q�[�:���:G�Rݾ���3Z�8��ވ�~�;Z'�Bd��J�Gd�|N��8�J���4�'k�r^ewN�o��Ʀ��e�?	�&�("�fUo0�a3V��t��X�R�k�@PM���f��V"�<��ώj�l$}�kW�ȹ,�v}��Ȋ�׭�+A�!��ݡ8Lշ��%ՕB<�^�-?��X8�-u�b$tR"�~��M�~���m�(CD��L�F���Ė�=��2ޝLn�G�j�:�uUs���>ƶ1���}��+�9T�g�����`y��
傁o�����cΩھ�:��B��de�}$���L��}HQe��I�wg�cg蚣2��l��=���j�_�y{��5���_� 	 p�m�x$�rD����zj����b��Q���f�.�9^+|Ҡ09޽����[䡃<�$6��
�|g���bۗ�!x��Y�kv<��U=O���N��hv�H�h����ZK��!B��m伴 v�'���C�y�"QP*���	R�)Y����t�>C2g��v��0�>��Yݞ��h�%+�����Z�Y�D.�K����>�s;�~!'�Ij�|����2B�u�h�����^��E�����XH�e�Ϣ��<{�N�.��L�*AzT\̲A��r��T�^[��=[�J���$>��{��������ʬ0C_wT�'�X�����1��t�Ջ1��@��U�*�Wu��p�ܥxF+̹���2r��ngk
�~=2xJ����b ��E�_O�H:����ڊ�~H���ٛԝ���.C�0�,��!�'�J2�	��k�t�b��z�~��_'�Dw
I��	�ȭC�+Jky�5G�~;1.>|~�:7���7_rmνq�@df�7}>-��5�^����N���|l�W�EY� +��ߙE�hs����4P���U�f`w�0������Z�.���i������ۦi���!K�\�{��wM��|����j�G~c04��_�����Eеhgi�5���	3T�B7�Vt?�P5 شq2�>���f��^.����ӕ�;����=1PY5�&�;�3T�	�$��'->��HL�q�7�`I�3S��8�*�fՌFv���+��=�lg|�
�9�d=zI��fa=��ڠ������@4?�s�]��<��Vpl��?t*�e�P�n�h�E+u� ��S#�{�/��,�ģ�՞ŉD�K�Z�U�E�W ��}�����;��^���Ҳ��R(��_.SNNk<�)V7<9�#R�4����	x�C^�Z3�Yg\��]���&:0�P�^��`���z�`߂�7�5�f��6v6|���>�ԝ$��ٻ[�N�(�`淪�:0����l�X99AR�A�U��7�lb���^���B<CL`� ��!���d��ȭ���EV���{�3^���ȁ���������� �a��$#�A��ks�����Pp�,6p��	M��t4�����tYo�{V��U4fkQ}ź_�9s�%��U.+�G�ne����@�8Ґ���dХ=��n:��"dJWUS���#F^����:��aku�
���\W�__���1�V>����(B�G����ѹ�Mb�%�� H/Av����]:k��V��㛫�gr#��8�ٯ�]�V��#�)Hh=��.-Vn[Mom�Yj`H?�3/(�3�0>��f�<�S��(�ڋ�l��M��ڗ�����1[ʮU��������� �� �`��ou���7�1[��4Qn�[��z0������Wa't�d��r�`��g,�~��9���MQ����q\�S]�C���꫘~��s�}P�9s �҈�%?'�����g�Zܘ�u�{����)��x:��j�2�y�R�2 B�QES?���&�5YXS����A)��3ru�E�<�6Y����GF�]X�:4�k�
��ȄA�'�J��[.R-D�:l�z��lʒ�����H�Ga�)����#ׁNX�Ϣw& �=ɐ�����C����  B���(���HS���(�g(�x�Ǻ9�T�SG \��e�D�=M��Ӧ2����9����t�TU��Mg�E����`o�$��T�}ݥ.��ǯ���d�rak�9G%����NnS)��Q���@���#(��L��f�?��o�?/�,(��<�,�9J�e���a(8
 �J3sT�{d����V%2���Y����+7hY&_'�oׯ1š�z�Ip�T�p3�S���C��\��p/�'b�ùl�,YA0  ��dk}#Qm���<����	+�	bc���6zS�D���pp@�n��f���Nb�H/����ܫ�ᐠ��C�̃��^��Q�JZ��Vz;��c�Y�xC�!�K�eKSa)�S�N�}h��;�P�T�������V�
�L~�\�X���f�a�]%��Ĥ|<p҅�Ri�7����R�$� �g>!.��N�DGM�h<R��%]�{�O��{��o�ΡƳ�s� ����W���dc[S���t�����L�u���1��rg�+�z�r�!u�CDe�J�ꦐ,�5��Xl�˥u�~U�G�@�����Y�;5R�iG^^i�l	x��9�MidIІ^���J>v6�p��Yrs�A���.b�rv�a㵆���c}���-�~k%�>��p��n�T�.WZI]ܢ���#�� [>F��U;�c���xᦥ.��~��o�n��x5����|�o|T�=����&o�x�12������-�O!.a�9+�%��˰���Q#t�fs�����Ȣmu|�wbT�ƿ�̼s�^|�-Ni{�����])`�9�J����! ��m�r{d��d�R�Ł�[�Z5/��(�*���2}_�&ǵ5�2 �sC�/�+�]���C� �
tc)���o����Jw������_a3�$��y�\�.?�!����X��`����� ���*3r1ez���M�a��,�YY��_�yre�4��'Ez]]3�����}�0�1�V��/�9]״�{��Ic���f�w	���}j�l�����/`�¬�#�,�0�x^��$sR�Q� ��	��λ��_��ko�m@Y��}��y�?��|lf��X��Zv7��y~��cA�M�n�8��Ko}`��	6�(K���?^�]L��}}Z�k�at�.���FSC��"��2�l��(^�	U�,@.7f��Z���,�G�d���V@�X`\�x�܍�~�o�C��ِ�i�p�;cw�	����5��H�P���0��`���E^H�(*���8��	�ߋ:��,蹒���7�+6�u�S��K�G����ߋS��dz�	����z�Q9�7`9sn��4���ce�(��gI�ZΝ-�VN��G\(�o�T8w-�"��1�zUj�W�V����"�Hx=�I!BcL��!X��P������ÙVg0��K}"��`{>�S���jW�fgi�Rяd`h����mxF�����Dc�N6�E�Y�<`��8Mw>�����)�l�N}$�\Z�ۡ����Ӈ3g�:��Z ���>����)]6�1�R��;��?	�N��ۜw�+�q��*8~Q�%9�x�����i�l��M�EgT���}5ھ2�؁]1���spml�{��\�����>"/���p`QՌ��d`K�M��I�i(���xu�XQ�@���H!���F�)�)�*i|q��7�QsI3�P�Y_8����ن����BJwp���.�[��q�sF������/V�>DaΚtra�lsad{��'��ܺ���7&`srDD'H��2v�{3�I�ߗ���t��&�]�"�.S�I��~�G������9�af�xX��Z���H���3���R���UV��D�z`bW�������Ԗ	KjXᒯ�Z���'��`Bs:)�c֘�Ż��\7�����84=4J�`�s���C)�[��Y��2�x�|@C��"P�=�]��<�w�}��;r��>S����0jh�+߆�e5�f�=�� +�&��{��T&iО�n'��5X�I�������ʚ�C�����f���Sxu\�9_ 	�!_ι=�������~*�҃s"�l��:V��Q`�.��� ����s(Lb�1�R۴Q���H7���}�`����H�L���kNHx~c�_]k5���I0Q��Ҳ`q��r����mi�D�l�媗Ĳ�� �鶮}P�މ5������z��u��p����]�ZZ����4	 M�7;cV�{u򒃅�n����5����98��!ܝ��p���?�U�� E�F��k��ؘ��
N:���P��	<�is{z��2ӗ�jZAR�j@o���� G��y��cV��K֊1�6�d�����9Q�&�b��7�Y�6~� p۫9""�)������,r���K��D�C��Q}�7FU�7�bQ�KS��xjy��	uxp�Κn��8�����y�h���tI����>ˬ�s�ኪ���l�Sr�㻽���y�����w"��L ��L@����ji�*�&����������EB��*c*_��P�=$xW�1�t�5����	aT�Q o�ʼ[(Yci��1�S�oD?��uTa��E�!F�H�6��Kr��4 P����G����F8{�~_�fd�o.�$`�E�W�##aA�~�ɝ-*�Դ��YT|�C���.�E����-����9�����/�wGY��9l���.�5�׭Cǚ���,Ɨ;�ih�lL8]OȊ)�1~�(� ����˓B�8�`B�v���Mܔc�Q��i�@�r�1�%	U!���?���:����]X��39h(e�݅"BRN�x9p3 X��B>��X�'[� �I-���ޱ��$)��j�>���Yie	s% ��������x�J<,@�q$t)C��q��9�/���0��v��]� �G�y�ท�se�a�Z�{TK�T�c}8��C1(�OX|`Q���Z$Q��	�T��d���|��K�e��G{��� 1�xѫh��G�#�3�'\7���X�D�ϒr���vI*C����۫H.A(��Q|yg{Q�vБ���֑��w�Jo�p�`y���ו� c�^���*D�� ��]�ž�E��2L�G�Ш�(�5�}�e0�Iw�#\�O�%�����+�������@ثP/oN��%�>�y�wL-Ö��;���T�$Z������)KT����I,��OcD}lv]3�����9jN�M���f!��-���(Y�]������
Q���Đa�+���0k�T3 �o�!o����hs���3d'������Mk��)q���aS��Ɨ�ۥ6�j�B-R�������2:���Z�:� �$��	�ݰdy,������s�9R&Z�����U�
Z�} s8Z��`4.����W��ՌZ<x�:M���p��E;�F.ҽ�ܼEو]��B(�a%**����@N{#�B�	��L��oDD�Z1��mU1w^��{��%|L	Z����1'H��B�������׵�H�D��B������i>�50{�"~�5(>	P��3��π�[x9����~��g��������t^KL�f�=_�=Oo<;���]��Z"%<|���jE��6*�im��R��T,*�����JC�yK����W�N[<�gz��M�׈�\7�m1:C-Ϸ�y$�-�lr��Ϗ��z��>y��]t;�0�ABG��`B6�Q�&l.�,��ybz�|AxQ/F�YE�O�;q=T�c[b �ɱ::�jȄ�,�OLM���P�鷿W���k}X�}����Z��渐\k��,l��qy����:�#����;���Ƌ�$��ޚd;���jR��~[~ź��E���E�e���X���|�|"QӜ���q�<6Y��rH��/+[�Y� $��ф'\�p��_g�,�~Y1`����k �//�a�H��ӿ��=����)*�ĵ���{�[S�s�PIsj>Xt�]PП>N�g6y�'K/��¶�5�!5�ߏ?�8ٽ���L���hj�Ԙ?��r��I5ڒ�j-������^��d�v|H�C0HJ�8:��aM�)Q�[U��[/{
���YJq�<�;3`�[�
]���KW���I���%^�a%l�O ���� ��O��͗�	�s]�$	�?�of+~�ٸ����l���M�Eʇ�`6��w.�J�5������aZ�A���� `��iсVt�^yo�ꂋ	֟�q>��MxV�w_�&3ܲViH����W���Y)�K�p"^�n	X}�=���L���ʪ�F�"=%+����Ә�~	����߀mx	Im������bJgd.�:�����66t��+'��OFJQ¹�g6�A� �����ϳ�4�@��؞�E�����f��?ǋk���cs���R��:@�A[�<Bgn+	���:2�|bh��8<�j�G�����/sڷ���I*��t�J�.��jȰ@�/_�����:#����?F�#n�����c����!��G۵��Y�F
��lؐVꅠ�-���zDYO첳C��V �u�dP.���c���R�ވPrcW�-r�05�X.{x�4)�e� r�#��e���Fۇʇ���f��o�#��D-�[{

���\�bW�4;H�:���aI~M�tI?Xg��%mh�����	껫��.3�	�xG��3�5����l3=���)�w^�oMq�ͽXL�ӨG�ڦ�/�P�E����5M`ԚL�u�_:�~mc���7L;�m��"��}��	-�5�P�#!��hS_���րKg����
�{���2�+n*���Ew��g@:>��cX����C^t*��G+$ǈ!���aU�b�Փ�S��L��.�I/��a��k`��KP��uOJ�ka��o"G�v��_��d��%K��������͎��l�u��SEq�6������=����3�(�4�Ux�]o+�cd�����Bj\�:e98�ga-�q��2�F���`"0czkEu$�
�����S�|"�]���Wb��&�Q�h�Y_���(�'n�3-�|��*��dZ���<v~0z�Iqٺ"Ew;�1�^��;�N�:}A�)��:8�S/����p�~U,aB�����X�.a���U�-|�  no+<qg�oޫ�æ���n��2p��h5���3V;\�T��a�?t�x�~��t����,㷋�����Hf��c���7ݘ���Lkqu��G����c9�h:��'�<��+{�z���k�$Ϋ�k����d)�Է��7�oc�Ѥ	�Ŝ9{2f0�Y�N�F��P2`��ANtAGq��sC�D�Rw�������R�]��`�X��2NNh���c�օy��<	��K%B w���m��l�x���l�d&M0�19����A���"_��Q/� F�2O��S
ڶ� *.�&YT�c!�L|TVI��&g&q��ٟ�L���T�L2�t쾉����v}��ԧ3�%{(G�Z�fsu�*�;��_6U7J�Sn�B �*����&�:o���t�W'0�7]$$��U�7�j?(�r����ơ��΢/o�6/��0��\�	����)�,��vw�g{Ē﷧��l_b�&6��+~u�Q�͜!��a#{�sSZLk��b�L�M�����U� ���_X�-����'����'s�o�܇ͽh]TpDɤ���M�Q���N<�X�W�[iI��9����[K�w^O����e��7��h��9��΀Ȝ�����D��Mu�:`Gذ��V����Z�"~88{��bg��t�?��-�֋�q�#���Aҙ0�l �����#�]�f��d��CH��1��+����~��U��gDL�3A��>�ʔRK����GN�ބ�0xўs��9k�C�����
��'���i�^~��-��Ax�����LP&i��,���t�}z8��B������������282�1rv��d@|=n�!A%�mR��ɖ��9o�$=!�_���P�)���[���j���~��.��gg���֚K���!۽�O�r���ۑL�=<���M퓍��ԋ�?G��_sr�_�P��u�g+��)��"G[�]�|p"�/6�k=�1�t	�)�A	�^2�����ci�����w�V|�'O���%��9�%�O�򽿄T�{Ë�1�K0/���P��uf	&�}�[��=MĕN��JTENK���"��(ѭB_�I/��-U�g�8����L����G�꣛-i�&g��iu�G�ὑ0���������ǐ�4	c���d *� �+�<������ �?��8��
�I�6��q�N+�۾�3䇊��K#����"B�O"7�<�M]��ĸ�aF�&��D
��X���H3�$���8�F{�A0Ԓ&�&_H�0	��6H�ި�Br=0�Iβ�~u��4݉��Đ�o�����������JH.���@����퓎m�Z9g��B߭d=FXa:����L0������_��	��N|OGc�i.ȯ{o﬒�d�T:'��:)��D�b��h��}�8�����a�6U�G��f Z��q�)i��^zl8Ƚխ]m�CIK`�2�&��t��D��-��ͦWU|�����z򦩞���tﭏ���|6x�4��w��u��v��K����ǿP�9f�<���o���qh�ǚ���� \��c�*ɺB�kQ ���+~.��=�b�������6(Y��`Qı�.ŵ�"k�?om��t7V�0�
�c�M%��w�+��O<�bƗ�L��N!{1�l��rm�f��\'���ܗj�����MJY���i�	�l*����f��_"�݁t�}\��q��"DA�g���5��4tf�K�A]b��t#��vHo�����E�Vj�&+�|��}O�r�4�A�v�gɯ$��Ngݿ��P_A�v�Oa���RМl~�7l�'j��?�Vn��ZTP��a�j؏��1�G���{] �I8~G�R��Z.������%Q�}�Xt�j��Z�`�D�dE5 MC\���U���N��� ����t-�+�n=���a�TRIH��yr�-���@p��b�f/V��	��$Ņ|��^zL$w��>��q��gu]��+�݆aK��%@)b���w?%������n���X�}��cl�}�Q3�����H����T��q(�a}��n]8������QAAޣ����g~���*ή�_$H��F��D�<��C_UP����Oy�y傯=Jf��`9>o��
n7��8E��>FB|�`��F,`���e.;ۣ8�&7�-@�΢�BH|q� fg����!rΙ�ݩT+�|&��)�&��q��9��}����Һ�k�Չ�n��S�f����&PM	�N�ZIՂ�-��Ò7��'�ܙ��#�P�}
Z����o�Q<#H�Wd�B�:0,E߈ٍ݄O_Uk��:�p�+�򅯈��'�Y�k��ނ�ޒ�{�Q���)C$�4`3(�u������z�]Y��JI�D���x.�q�'�c��Fp=��
OΗ���������gB�ؑ�8�����wZ�,h���s/�Xy4=U�N4�g����g��O �Xb�
�?Ӻ��5m���Ze��5F1`��hA�w5@[q1���/��T��)�����?�ئ/��],��i��� #����T|�h�¸�%�?fN(��@-� .��Z� �h��1Ƚ��qZeg>J��n~*�h���Z�c�x�<�F�8�R&)[�usd��^�|���3���+uN"��[#P�������������� ����]�8�*��Ke���`�	�wBR,ܤ琟���v�,��(�P۟����m����i)�%�Ml�Ç�3�ѻل�Y�dk�[�6ꎚD���Ey����60t{�����������4%�(��1u�ʬ��B��x`��-�rn��3k?!�,�2}5J0��OB����B}'☫F��k8����.+�&������܂��X�a��l�oU��A3Xy�szd\6������0od��*1j�g�-j��0b��Đ�C�]�U����c^�߰fY���9���@�!�uEPW��� ׫�Y0��I�髏��p����%����no1�.l��Y�٢���v��6Apf��D�sZ`�O�I�4,;���'�y�yed�]4��������� S��� m���P�~����Ή�=Hd�6u��d%�T��v�����z)u�D��>�8�F	��
t�BKMX�41¶�؂P���~�w�7��a�ooW*��ƁV�M���4�X�A�9�@�qd]ռݢ��
 G1p��d%��6F��7�K|tQ�)�H���)���]��5 �p� L�*��2&�����V��t���e�I��_��.\���k�"Y ��'��\M5
�R����Y�f<536���0��B�����M�<Q��h��#�9ՇÜ(;�[��.�g2�#��3�_�A��q�Bm���R�)_�wkN��J�#i�k+�Ӫ��=���'HgY9;ڄ #Et��!\�7vd�Ԅ�N���-;�Hq�Nr��x��vŃɁ����3�K^{d+.@4b[)XS����X��E���&&�g�.��r*��	�Y��Y�4l�L!ҦVw.�f��D6�T:�r=�r(���*��D���,2��Cf��
����*@�1h�� G�q�xX���	���Rn���}���b�t��x!�]���[��Ma�,�Wv�A7<�����e"�P> ̪�4�cO��5ɛ�.y^�OM����K�9/���A�@<5�:N\��9�Z�������-�4�C�p��z��ј(1u�e�O'���Ƹ(�Z$�~� �k���'%Eލ�o��Ы�֝߄�UM.�9u;H﬿���e��U����*R��W�7ǡلD��#ưv�9Ş��p�ъU.��V����iA��R�u@��1�k)��mp��X7DV�?�J���h�öN�<�K+'>�y�+���h��y*o�V��OD���H����3�=������w��{�J��fr���n^�MMw�9F��]5z.Wޛ��IV���~�0�@��X7p71�g��Q���/��=�(����=ox�/�d����H,�0��tl��~!*V���}m�p�.��e��(�UVy��F�����ȥ:�$��rTҷ��G#d����s��}T1��,Ə���g%D-]p�$�?$hn�U�E�k��fϔIs�u���%�#\�<���\��֙�=6���Ѩ���dA�,<ˋ#�Cl6�w2+��Q>�揄��"�٘r
X>�	.f5ڨ0e��#�!2������Y�1>�#}���%��Ǭ���5�RT�j�+�w���F�Pj&���]ܙ8��e//�T^m��{����k����_x�N����wc�,�Gxy��A�2mC*w�E@Is��o<a5U)�<�BKArKE��6Y����)��������{�#����D@'��n1���;]7�CR�\B����[jr�bW���%`�H��=hԶ�m�uZ����(��dR�3^ўJQwS+�+�5��<k-�K�
$;F�I(��5?YS)�
���:�]���8z$VR�6F�}��*L.����nN��Fh�W<�=�����'��]��}���7��l��io��Z����C$ ��Y z^��}5�b����2}��v�ן5Zo
�kl��H`ʉ�`������}���ɇ�ML�	�[�qB���+j]a�.p�
�-m˭�)Q�#��?(=jB@;��N�2�8�Ϗ6�Gk�q��ڎv�@����Pq��ꀫL����4t8*\k�呆�R�>3�n��|$~$��*��Z�,n2�aћ��^G�;8�\*Qe��^�q�����7�b�-j�%E���4���@������5KT���\O����V$�,�����F�Zxu�J�	K4�ֈ��ஹ7��(���R�Bff�"wB�W�j�; �sE�3���`�l�s O�̕�i����S-�1��a̨s$IDj]�ל���Gm�d�9�Ϟ��C~0� ��o��:FI�ڶJ2.��!4��+K���\�H�Z?#	� "Hg$�ss�?����~��tO�Ɲ>���#�����\��ұZ�-Rd{��������~�\p诋��,�uq�sn���2p����8�1J�6p��S�����n=-x��aاd\�Blu{fk�q�ޙ
bx�OxA�j�A�e����0�᚝_2}��/V!B���6�J�9�E�y��'��	'���6׮�5�R	�4�ԅ��Id��۩yz����m>��r���?��b�����u�U�@��䢂�Is��$UD�|��FY�e �V�Q��<۷�PX�������arE�!J�Q�����Z��K��_��<S�N�Y���Hq��YN��r�΍�m��8O�ix�e麣 ������)'}[���Ȳ�z��*�s_T%9z�x��� �t�ژ!�Ց�zS8�v�m�
.�n���v�S�_P
��<�gEӦ�:����Ԁ0K��ǻS`C 2H&�.��AZOtMa���4��K�B�<�FV[��r*��B�� ���LQ^��(�5�w��TD�"?�Vn��'��VA/����+�����T�7�?.���@J�Du��>-���yw���+."(�3�C�0 vNt�[��VP�4]"�D�N�Y�(��Z������o'�-3�S��}����=�˙̒ z	z�r��%�$��P�c���\9<z�f�I� �g�_ ���4��\��N�ߧ�k�h�����3ˇx�����Nlve%�P%5�Y)�x�O>�(`�|)�Q�6ҭ�gO�a�%٥H�s�D]��QUJu�a�~�a
����^2/����(tK+��E�h�=L�#MV#Z����q�o�o4'z���L'�و��ٴU"89�����m#�W����¾�F�����N�6�hX�_ J��bT���Ҟ�µ��Xj�r=9���rh�}�A�r~<V��*$X�@�������|<E(��W�D�]�m�:�rH��&G�����^�W���Т���/�ӊK��Y���"�Ȣ��b梽�Y]�;�!O�KQo�����W����0_)"t����o�VBσNĒ����
eX$s?�P#�5��K�ɫ��	�e��g�_�i���k+����x3�-�L��x'ל���^ �s&u�u�~.MApW�&&e�ՙ0`Q"_�CB���<]`���3P/:�����@2���`���|�$j9�r� �>�"��!��ʈ�_p�ʤY�\#�/y}��]{z�B�]�JC`܄Q��Ή))De�!��< #�9��2tM�C�DDr���5���w�j���+3r,鵂�=���m$��֎ c x.o�Q� �,��N��'��+,-<��vk_@}:Ɲs0kԈ�/�e�3DrT��'W�SK�o4&�i��H��O\�y�C�PM?�,�f�>� }*���Ew)�M��G�����b����|d{@��\��9r�'ď5;;���g���l�.�n�@�N��ך��܎%A��S�uˣb
��P��*���.7����9^�-љ�T0Z���0�¡��<�����Q��&��S,͉�kK�n���\z����E*K�����G�����N+�]��3��b�m��Q)�Ŧ9�9��1&�Y�0���;�*�ڟ(Y�n�ۂp0(�[C�a��,���o����U��U)$4V�����EC�5G3��[��}"�W<iG�oR`�?��l>�����^tx�]h�a�`��<H1���`H2dal�ц�U�:1|��]ll�#�x�:蟄�5�Vc:�n�A���B���؇w�
�#gi+���-��!η끆/wP��i�I�>"�u5�E��B�5������P���b:��S�M}�7Ʉ`>�5����h{���d��Bki�}�-�+�2!��6�/�إ�&�%qr�o�Y*�2���In/g~ ���Q��M>��
:�z��ʕ��0��3/���H%<��*���^F"���*?����Q��:��f��^���P�=\��0pQ��bt����C�,���b�9R��2���6J�qj�&�q�V��Kƃ��R�.CY)@�F�[cH��2h��e��,����q�N��9���x���n�D)�Х���wF�d��Y���v������݀���_A=�/<	X����*�a����_(ysb��2��~�- _�oA�*�cR���>%�7�2����J�LKmԖ�T��53o�����)����ӾWԗ�E��I|�M����ὣ�n�|G�
�P���������cBϮ���(ï�Yu�ܨ��Sg�X][���^��F@�勸�I�]���0+Q�-�֙��ߨ��tW=��h5$�;�>�7��{��^�#=)�J8�*�XE6G0ic��*����\B�{hXjf]Qp_�m"&���C���)�wT��J�S�5�7����-�����R��_�IXڨ�Eiuu������	��s������#YT���,�":�l\��^Qy��C]QC0�S-���/��#�j�)�ATu�=}:f�U#u����^oQO�{� 0�Vͤâ$a	��IrbOϑ25�
*/6i��b��Q�@�0��_�9��0�c�j������T���� ��ܫFn<�a�Ч5P�Vl���f~����3��T�&2˂���z�O��)N`4��W� �{���������f�펄�6!�P{�_�F�ys�k�|^�0�� �Gr�[�dG��+�N��_������_�SD���\>�K�`��R�,����� r��x�f�0ȅ�xq�h�*�&��h#���[&D<QU<'
=Nd-G�����ڴ�xM�Fn�#�B%��0g��@�v�ڪm�N<&;W����_-�8�ș��<�8�O1��D���oΙtCj��@�]�m9�^��"�J���P���|�����\�Q|�0 ֖%*�6�g��H�#.{�PE0��<���o���+\���9t�����괾�q�qxO��-k��s�rnv�ܤ���1k�3I���)���eAJ�5�P:�U{ ,p#pxA�urU&���e�?/�#��3�aٿVC���]�޹(o�%
��eE{hS߇˗wtmTEL��{-�}&��Ū��-̓SR�<0K�:���<�#M�k�g���z�
�k#:���)nBFL��C��Mc!�4�4S��N֎gin���w`�j�5���Xp�=V�mӈ/�Pkg�o�LԆ�?o��ə��
B^Q������n�q�G��lӄ�,L�C��ܤ��0�P���z.i���,�I���f���X0Z��籓Tl���Z�(���l[fZP�CXY���l�
\��(b\b~��"d���Y-���b35�QڧZ榤v���.���Y/;�bِpx��y�����cGG�I?-}gR�a!�k�Ͳ��1e�F��^�!�.���Z\cv���,��fT���^�cW�=W(�^�rX��:�v�l�
 �� P����4⵵�P%ѧ���O?Q����p�`?��=xTdA�ݲ���Od�Z0(|	R�+~�
��E�l�[-�\9ʺ.�>K�F���@�,�@��]�� � �+j}5B׀�# �m7��R��L]�F�ŢE0<V:����x�~�S��� 	@��R��<�)`�*z��`�pG.�
��;O��Ǎ=^�Q�)B'�Z��h� �Qí5�Y����o=�[�уCm�-'��gyG1�qE�#����4�2���l��m?O�sjX?.k��
(/��+�t?~�)f{�.A!�e	ecX׵C{���i˴�M��seŠy�v�H���rEr�{l�$z�=rLZ���@cy�Cb��NR�6�нْC �����z�֜�0}������c�{ґ	j&�x&�쵈�|�� &�0\���d�Q�ϐ��`�!�4����9��}��g�Eb��,48����N���ܶ�6��-���Ǥyg?��-�0cޯ�0�7J1>�J^)���ESu��j�S����]��K�=��X� �B�����Ų��=�����e0�����{�F�I�� m�s1��¦���`ε�Iȇ�m��!�h�qK<�>t`�N���y84�,Tׅ���!C��w��Ap�GA�(��u+K��-V��0�5j�1��`,�=���n^!�/���r�E_��Қ5lP9�5��{�~v�<��&�םj�3�,U��ǟ��֡�"rg�����Da=���g}g��IUQT9��=�p�;&!��JK�Wx�o���tA���ԠJ�5��mV�]��FVF�L4I�4��qliP}����4Ҝ5o�1�e�����t^�ațߦ�,�r��� 2Y��������C�m:մ����n�E��L�xM�!������Fj�5v�[$-��-'P8������ ~s@T"1���$�b�|��J�!�$��:����g�i~�>w�tkW��_���w��<�A;:���w�o	��e�p><�5���RA��yg��iV��-Օ~4 �g��|�����|8|*ҟB<�