��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_�}ܛ��.��i�F~�~{�J��C�a��K-?�<�>y���yewY�&�_��wr��� jK���w��C�Hxj� ۞�
P�D
��6⼞-E!F8��ؤ�Ct"�<&8t2%A��G9ц�F1�#Zl8���<P-�J��E��_i�y�$=>y��o�}籅i�n.���%c�Īѿ�P�T�]z��U�XpQ:_c�.6�]%`nK%E�ijlV.5�Aa��������x�쾔��傮f��+���䏦�P9���o!�F/F|EF��IkՍ��ApD?���9ߢ��o�n}�����=��O����)�C6��m૊C`�<�aV3d�;��j]��.�L�'uϽ2�d~�/�1���<�n�H��x\'GmX�y�`���w�6��!6���k�l')���)B����A�9=�T���ڢ����j������_�\��vW9��vuF yP���|,稽�f�o"�]BeN��?��n{�o��ۥ�
~�x\���O0j{�B�J*.�.���8�Iʠl���� )�eŔ^S����w�X��C��F��q��E!�˶1���\���>���j�3 f�S5���^b�G҈Ik��}�ָ�6ߕ7���F�\\up
��A��$I�4{���n�|�4�C= ���c-�C�ZW������B �^��S���Wy吆 �e�bw�6a���3���U	)I���9�$�"��s�S<VB8��!������S6���܍kY/��%VB��3�z�>A��h�2h�ܠom��a�q�>��[��!#��=�,���f+0�Ƽ���@+#@����W�ݘ���,_�&�U��(�BS��ʈ�����'���1�2�5���nZ����ڜw;�vL�^��w�;���/�� p�)>��� Kyw�`��é���D���W�m՟v�h��s�&[A�)����W���&)�#��g�`���'��%�������&S��2`K�^ޡG�-�	,��h���6�F�#���y  nB��}���M��Ol�T��1���� �؃�v����#BtWn�#q8��ώW`���)\�BLbۑqߖ�A`�[-�����!�ZI7�^��X�Cݕ��7]��NBU�;z�W�ɡ�1����I�9���]9��f��Zc�- >�NbȮ�m��?�d��MP�n>k�՝*���y�.^�w�%*����՛�s.��ԗ���Ffd}����O�LFnP�s!���7Ǹ|�amK[e�C��CuL�$s�?��iG���w7�>���i�P��  �������BG8
�{Y�L_ ��|����@����l��iv��Z�>��"�|A����Q�+�>V�ҩ����TB�8����m�/�T��ɠ���)R��t���<�b��X	��-hwEo/�=vQ�{�-p�k�x�E��e[�(�/}CYHP���}��e8	�!�M����͝?K�n?y����yssV�Mo͂��~!	t5�^���C�)��3	�	أّ<�v�G����l^��ϖ䙓-А۬��G������v,�p�!0<0{h�V�}�ɽ�ų��~�Xn(D�r�H�	}����6;!+XȆe���xA �J0�IL��Wt+i���gmrr3��@vZ�$��8`���6�Th�#�✾,���%9��u��]kڸ�#�vE���A��9a|T%�.�|�c��
���u�sF�p��M�N��|�`�\@ )$P�����ЄGctb��]�z��4sP�)~���U�)��U�x�̷%劁�Υ���e�����q����sOfQ�e{�5`��.�`��c)�c1��=&�����y�T�װ�Ni3��f^��}Wo�-!���k���q�?R{A�׋�U�D�yԂ�����;]���zT�[D�/���ͽ���g�4Px0�Tƺ@㦫�B�zfQ�`��P���w�z�����@��۰~+�|�Bm�3Z��ݞ�9{�y�̥�t�,���He^�^js�p��-%#(=J|H�?8^�{o*5����l��t��0U�7�|��|O9�c7���).S��>c�ߘ���B|;�o�r?�CoP[�,�-��t귛�L�D���$�n4m��eS��K%~��]Y���6u�������6�I��1O@��-`�,ޣ�7eCa9Vn0U5p���,�G�dcN�t�h�{��5g ��� ��6�lC�;.��)�/�u-�v�cn�V������vLmqGHj^Ŷ{߮ϡ���6Q|ܳ�>t����!��[���R����f���	Al�|�q�s���ޠubx?�T�Њ&7g�����#�G.��/���ȃ����pyD�9q�{)��e��Ù.�D�İ���]4�@�mί�F@��T`ê���6�V3�LS�_H�b4ϓ|��W�s�Șc����o��L.��&j�/ï������������r�$]*	���U�ɬ�=�2F��(d`�+�_	�9GY����<�6��f|�8-���ػ�r֩;<K�K��v#�\��¤���S�Cf�xZ�"Z�e�����å��2X]_Su��06�������۹��!ɻ���Oq!Abm3��M��D�x+4�!q��p��yl���y��4���ۗWZG�l�/:%"39[�jG_���y!
,�B���k`V�� �BO��_"rܽײ��mY�gr"k7���`�N�����&Q��kR���z�?wcq�9e���w�v^��(�|�J�d�>���Qo;�[�����c&���f�����]q����ޓ�v_DV��~5�Q��9�ϟc���KSi���Ĝ�ﳅQq����g�0)�� ����-+��)��gډ~s�S����7gP��S"{I���|�Q�z��!޶cKD��t��-�� �,H׉���^�q�4��yLf��unn��/��g�&m���r%�RZ �S�u��W�֦?��"�y�]?��d�3!�ޥ��`�r.U���dgѷx�o�?8��'6|��t�=��M�}��U+3���h��	�?�z��|fo����#5��و��/����_˧�	�����%�?y$�c�.�o:˘���k��Y��3�/#�0���:���0�q�X� x������B�l�bc_��6��\#��tL�=�!A��b'2��J�Έ���O>+�t4 i.
�>��H.*HQ�?O@��[�GPN�Y(�y�j.�|c���f�YsQeV���/������5��Q�S���8����/�1�3\1����H5缔�6`�f�e�C�{�8YB��-�,{0�v6������`�V�(�W�k�n�@�_����N}¼ ��-�l���5v (CC-�++��EY��a�5\�|U��ן��RWg.���;�5��_���z��ݶh�51�K�6�=>K(�s���bRVq����>�;ķ��ȇt�O�6�@���r���q	��s�����88N����*6��X�:ZC}�zSa?R��8RS	�}d��r������\��[h���l����+9	��*_Taf?����jr�d�&�� ��;1�$�����R���\n�%CI�$�M^��H���w�����r%�&[�/��n+�kvX"~r���
�IcZ�-	5�W;�C��Z��`5��aVLh��K=�㓑�Vle���T8*��� �4�*1�l/^a���k�ݡ��b���(F�9�&ϲڄ{�^e����m�j+B��)ϕq��Ym;���|!������8n�?�20���fk�^��״���&�XEp�7ԑ����~�t�q�hw�J-:�yjU�5R�w.��ŝ�d{䵩Fk�"J$�+�3k(���x��1�ذ�qq��u�J���E;�>Y�=�B��ǡ��Q�e�3�Y�L�*�9/�1h��V�SL�n��@ӷ_���.BxL2׺JiA�``"��	͎���(�x��Z����B!�/'�,fd��r(V�ki��S���oyh�
�;�4ݴh�:+.�%�R;�R�����ֽ:��vwA$�h�͇����f>O�)/B�d"�vH��J<:<��иINf��k���|k���t���O���6g�S�~��*�����$����-����r�6�B9�����E;_x��`��W����Ή��|\J^d�[K:�q7 �q�_}V�,'���q�Us�%sVT�6G���bJ�&�D����y���+���L�����v��	�IP�+bG�X	0���aEj�U�aM��Z^B�4R������� :��1��m�Z��O�R��NW�M�w!�4��eW�隧,U�s|Q�=E�~M�*�V�Y�T��,���������X�y�q������<Ǎm�UWWˤ%˅�W��jd�X��p�q	��U��[
��Y���yhg:�^m�ߗP�;�'�����M?�s����OKQ��̰���H���4�/7������{7{�9$��>���t{�QdC�R�I��H��b����o���u�v�X'N�}� z4�M+8�*��tI�0 �!ihij�2*��� ���*(���~��[Sj�9ZH���j��ku�Pug&�ێc�ˎ�gu<E��3�
qb��ʂ�R�����31ɱ�l��P��3u���8乢��f04�{M�������1�N�-]R�g�Nz�1��E���i����"O��5Q9�^ޒ�������d`܍ی��o/���&"��>䔨�M�C���_K�[3*ShKSܬ�WhM��Q���Î��8�@����с��%v��.��=
{zw��+6z���yh��T�a?'R=�oX��0R�|�%�Q	^�m�z�k���d��OI�[�)��1�"�w>h������w:W�Õ�݉���4x,}�GO;��S�7��\�SiK�eڂoN�,�*\h��<�8���iS�A&H�_[X�mf�����v��X'6��K��E]y���A�fM�s·�����*���7�-V+�W��Byx�/&��M�����H)���h��JN)5�	�l����� !�;+̆r�M�r�j�mjU�n�v}&��л��ID�O�Q�*f^gi�h��WK�-`��[Y�-U�AKR����6�X;n�ݝ��0ƹ-�hk-��X��#���HP��p9��J�@�G�3[�[��X�pj�
������������ĠX.����H�C��׀w!L �}��-s�_!\� �9+e�{_@�Eύ��]4MV�N�(���K���}�F�؎��%�����I�i�C����Y��̘�:�?B6��Z,�����&�������?'n�t{�ү�M7����h?���b���Ծ_i���?@-}o����͏/8�!��$fH//g��h�K6����3E�^��_�.��K]�Z�X��b!z��a�B>s��S
�	ɳe4&��Up���O
f���m���������By48�n�ƭ�4�7���܅�S4%�h\zM��٧ζ�N��F��9g���KnO͕��k���$��CE�ҽ-Y�]�BB^!`��Ȗw���#ƶ����nU��w蜖�2�Bp+!T<8�eA�%؆��a��߻T��w^�E��ӛX7Ȋ�܉��*nD�A:/I���C ��U1yo���FW���|혿rޮ4��B�7�2��F�`�7ωPL��H?���<��Q�ϻ��,H��ǭE�)"0c��_����'�ةȢ;��i��
�Y�1t�Ļ��޲�1;�ժI��R�m�~��y#ua�5�	Η�px�/�Gmئ�[0�tܩ�	��đ��Hћ�*� ?Q�0��v��uf��3�о�Y��o��x�^�r�)A:���~mx����6�q��+��ҝ��F!r��6'{(ܗ@%����WO���ݾR�6c
��j�;\+�6v#�4�/�+1��|y�'�ٌ�`Lz�W�tTB7��|?VF6�Z��1�b����.��*j�8$5���k�;�P�L�5��aN���9G�h��~�P�}����i�Y�L����f7xe0f�(��$��()I�W a�����iH-C��Oxl���mU�+��z�y�*�_ܒ�������� hK�������|�����(�Ƥ��jt�jw
���)�;����}�s��Y5�.�p
������9�
����,KR$��Me.U6����q'0����ȆJ�vzN�3@DH�1����]���97DIGw0k���0��:�|}�]�fǘ�����fY1��A�@!ڽ�����c�O;H|��֤�I�㡠a%tS%lo�������Q�2RD�>��Qĭ�#ob�����7ͮ��J�}t�.)=�a{?h/���j$�g��-�;c�৲N�CK���hfYcK�F=��I�v���Z��[V�;D�����R�haDUq��L���d��(.��T	���nh��bA'ܩ��/((�p=���VŌ��Zƕ1$-�6����
��j�塯3�$4
�L����$�ms��h����I­D n���]\敟��f��j&p�-��ǲ#D ������ҙ���;�'�p�Ff�.�W:M���<#in[��`�� 5��]%�
���pR����'��"�"�P�b]�*s	�ze�k1�����ɓ�c���j�m�{l�"�Z�I��epBIrl���V���m�$Q���f�����8#+�@qe���)��7�O����Ӗ=�F�����٩�]#�ʖ�/�.�}����#��(9�R�]�5��O�(�eಕ�I�(vDm��:�.]߀|;���I �|3D��i�mE>h?���aS�o�LF����tÎ� �5�G�H��h�Ѝ#�kOUе�Cp�4(�z~�b�=V�ɻ�b�I:�6��7���.�"fe���Еl������N�M�B�>׵����p�>��;�O�E��r$Q�F���`X�Q$�ILn�0�3��+�CM/w�9��FS�$47������'%�2��� {\�êyNH��8u^�\l�Ր��ƈ�U�Ce;)����z�\s�,p;�d<�I��Q��K�pOi�6C���U��,��24˓6��LV(i`����Vu�h�c��e?��N:�)]t�{u�dR*�{�i�l��-��*�N$e�ʤ��o�U� ��R1��R��j~z�������.h;C=��c�����Ӫ��������3�f�\w�]����Z�ww5'
�w�����3&�FR2d�A�o� �n%�z�aE|�o��=b��;�J��@A��1��g�m�	�|�9�w��d��P �i�ј厌��^�\\��3$���/�ޓ@�����ٵW�,�.���e|�Ux�U�<m�=f�{�f�[���h�Hwl��?K{q�����O��,Dc+��O��ۃ��ӊ,�f ��6�MmAcM�_��Е�O�x�K��{��ǜ��M²�ns \ Nrv�� �����!#��vP@��pJ�BQ��S�'���q��G�ʀ٣P��G�������u'e5TIm<�`��f���06C��rt�b�?�ߺIAIy��.���ؤ��Kw���*_d����S��\E�Y�(�˸/��.�z��D����+D�l���@w.��`�1�e�q�_3{+A�S`�q&P9E�A�ӣ��n�N}�f^6�;_���!ȫ�^�O(z��^��ՎB��^_�Q��ذ��1��ᎄ
\�$��B|�1����j��u��S�	�������&Lq�9�:���j4� c��T�-��e�4��6����4�ʅ\�RAƃgA2vje�,߯]jCWV�����9͝.U�<�2I:?��7��ѵB�w�|5L������+N��@������ũ��uO��	S������ɱ�A��h�%{u�0"ݰ��X�����z�z��c��f�Hbw�"��mbfX���y�C%��~�%,�1�mյ�2�����ĩ:�����,�y����_�d�_�ۑ!�>�*�	���������-�y�p��f��������*��D����0�d���MH"���^���/F�B�R�5��I�u6kF��
�ak/��
�� �*�Atxz8�;�x��zH�m�Tݵi-n�L���H��z�ЄN��Y.�#�����KL���1_�B3?FS7eg<
(�ȻlS|�a@\?�L��kK� �������)�8�.m'� v[	���vǪy������O�k��N,XF����\�l� �����&Ha ��^{ ��W`c�f˦�L�����t_�z��|�͆�_�{>�XG8'��'ϸc)��G����ﮞ�ӂ�/I�	�Oj@1a7���� ����s1��F/4!gCu���p*(�]��&.�.�j7\[�<5Y@�^����n;�ʽ3�r�ۏ�w��7�?̨��w��z����=�oy��/��Z�Z����h��{ے^T>ۅ�h���������rma�@�͓�t���2^�q�)�{W4n|�t.H�h`����[-��a*�l�K=���n#������/!�uzJ�eM���G�m���\�tm�M(��.	p�U��D�-�`=X�.�^�dI�J�3(��Qnw/ �B�ҫY�nP�V����%ݚ����&��^��DM�eP�B���Pw���������$DO�͊�lFUd���C*N͡��NzacQ.e����ZV)\a;�+�ټw M��i�Sڹ��Wղ���?H�N$6W��.]��1.�������4�P��!EV؟
!�i���rp	l(�nʺ	4D���+���c��7j�v�n���7��r�2N�W��=a΂b�W��Ϭ��Z}e�ϭ��.���󨵊���)/����ę��>�B~pVƓ��4԰���3d�(����MG��˱8�
@��B���0��NO��8�H��ʻ+�E�;u�T�����[��C�����(^�6Z$���_J8���&̈́]1��ߍ�=6C��]�E4��K߅|%O�Wb��T�61%
�?qW��&�r�8�Jd�x�#��"��%w%��^���P$���d�S��+�3a�1m�\����t�B�&p{o���|Q��K��Q7�`��.����ې�뿐��>�t��䚥PU�d8<+	7�H(?��I�l� *g��W	��b���Q�ȍ���Hz�yX����^zY�hO�����ᓏnQG��G�: Ց���ʒ�,Q=X�7$eX�c*t���q�i6<Όu�;pQ�`|���?����;�P�q��r QD#J���pV7&5w����5���3��f��׷�F.r�����a���S������l��9ަGD.�[Dws�$me�}��0���_���;���(Y�����˓XhE
syP6�����-Â��TCu��ڭ��[�u�,���4;E�sN�coX{w�g�f��;*
c<C��̪<@j�1����y�E>*�g @��fx���lW�P�T�YJ��^۸+�z_�k5�f�4�QLT%s����|���Y2K���0�}����F=<���ygB{���1��ԋ"f�ba��z�`J?��������+Te�0/��H��:��ӂs�a��Q�a������o|κ�<q�	�;c�B�w\�����&]�Ȣu,�g�B��]�d��_��"9c[�߯�Lw�Ȁ�5P��e!�����G�ѓ�߲_]��h%�B�*ߤJ��Q�F�н�d#��!GS��,��c ��#�z�t��7��ƥWiAЦ�l�))�rd�vo�.��+�
��f��͇�7Z�r����{g&Ͷ.F�A`^Z𽙾���IJ������Wa*�9z�g��W#f9`��r��G��ɿ�8S���p���#�@aշ�����;N���UV04�ݛ6mN��Pq��h�k� ��Sq�}�ւF��R���8r6x
Y��'H�p
@̶��`�HY�Sgjf�
܀��R����Nq)��8��sW��*z�v�-r��"�O�Sx'"Pc��v�er�.��f&i�(A�;L���9m���o��_,(9f�fTΒ(_�=e�M�������kU�^�- x����{�����`Ϙ��K�7T���I�F�/�#
!�Z����E��7�����:v
�]Z��%b�E�th��������L��jSe���}�irbR�3P�8ab���ҴyD�I�fͫ�\�n��>p���L�|X0O�3�V���9��@��0���{.�T��I�W7>f���4��P�E�_��{��:C;i�;��Z�����.Bl�����A��;�ҫF������x¯�D-S��9?s�m�$���N�7����sF�,Ob�7���EB�~���{�㿸 ���x/`�[���� �ξ�3ɢQ�*?�J,��Q���z�y&Q<���!�`E̱�!ޑIM���F�?�&LC�R=�>�f��`����d,�Nh!��3��L
�ᨒ�b�a r������#�ä�{���)�'=���\8�����K^x���Z��'�1-�eZu!�C�U�2��=����E��X?Fs�K��*DT�l��]��ӎ��D�c�;p�^F64(��7K��FiQ��흻�EGb �15,�	t��4� g�ͨJ�X��S�+��.l�6(�F�e��7��,�bk qŠ?���E?p��A�P[�g�CUF Ԕs�͠A?F���,݉��1b��,�3��ݮ�-�DZ������X�c���TB����((D1~�5�Þ�~kxH�yO����F�@�Y-�2]�,��gFB����C8(/\׽{�B���ˡ�T�o��4��V���M�g6v��ar15А��hB�IѥX�0�J�9�!��!C�.�[�_��0R���od��ܯ2�ɏ6~g`m\Y��R@�+�-0�G���d
g��Z�!l���X��Wb,1��)r�X �����4v��S�?��W.Ԥ�q�8����$�6c���u6'��V���y]�͕����:6V~#�QC�a�W�@w�s��[��q%��|c��C?�a�R��u!r�,�b�CI���/>6���_yC	y��~f�j7C�x8�E3� ��Z=k%��� f��5L��m�W�j/K��S$l�^�?]xle�4ѿ��Ȉ3"U.�w *1�.!A�b���n�~�k�B%/N��d��p�h3��v�D�5|E���Ⱦ�@q��'���v�g�" 9��n��������E��-�T ��]D�����]��|�^�b>�f��5�£C7��&�{5��n��~c ���7�(U���	��K���1=t�T4�$9K戔$��O�$��|�������]����T�<< �J���[O�;ܴ=����&)� �������w�x�֤����J�(
����_�6�Ą��x9��ߊը��$R��y��@�By{����r�X���,T��YZ[)�e��E �M_&�4�Z���1��ќ�C�q=���Ƿt�U��[9�6��$���Hʚ�-����R���C'Wa(!wg���"l}�l<�"���X��ω��?{o��O~�^�Y��O�֑&��	-��*���9�ۥ��9"�dJ����6\8��m�xL�"��c¯�����|����<eΒ}6���i�D:fJ��ݤ��	��4�譤}f���nbo^�<{�K��>�����ud�g���l
N �Y�XPm��Vf��)���`i���H��5x)�NØik�����J�yH�Kc�@�ۗ���������|�� ��� CZ Y�2���p�Q�s����F�J_�*-�xzU�)Z��5`S��H�uL��0[;�<e���r�A�@��u���_=�ws���VRe֩�ͽ��Wʅ�+�[�oOZ4���xO�6a�:���9@�e@~�K���"���O�P����NJh�x�a�\JW�آ|����޲Z.�S�7o9��rz�k�� �I�7�!�G� ���-�î��3�`����~L��5hfh:p��:T��h�BM�"p[Oo�FH�Z8�H�RD����MR$��S*������A����YUۊ�p��P�T}�@h�&�~����
9c�c%��ŝ��I	!$����`M�v��Ԟ����Y���	Ϭٻ#&קE�a�]Xol*%A���*�hQ{+�7D�jW�Rp�]���>���Œ�;Ї�w.*�;���>wlv��b�Hp��V{�p��[˚Y��J�p�H ��vO:���Q<���]V�=c�6PU�?6�	�Q.��	��b�~��P�f�t�(�E����� ����'�M?�����71���'�=�kư�N�n<@>���xDFj�OW�,�S�΄L�n?e5PȂ�U�t�_}�6���?J`Dٌ#�=: ��@%X��TSU7*�-�)�"�������d����sbm��X�FZtS-#ؖa���Qw��G�%j2ZAY��=�"+;"Q���P#�i;�z�	UJ�6A��0坆���`��d�B�b`$U5<%��1zBv@!�Y3E̶�9�C��6�G�Q�(hP݊4胄�����1�\@Z8����+N�����2�[&9�m�`���
(�f֠�չpi�g��y���Xr��T<�#=���޾�d�
�tDp'8v�fg���ʖ�*��ܼ���@=�ۈ��\�2�F��}�~�v.p�.��l�UO��0cE�t�p�-��u�@�'��'{k	b��#ҲA�7��S�$�c���y��/���gc��2T�V�DO�R_r�������n c�`��dlb:tB+M������ҥ/�ϴ�E\��v	4t��ja�n���PE���4��Gp�%�pGoJ�C��D�ˈ�)*σ�c�}�C3���B	�&	�vBx��kN�o��.����Ed�.%N�P���!8�|��o��_*��7nz}��,����4��Y23^�%"o	o٪f,�[m���'Ƀ1�`�����)�ܭ�Yx�Yb�e���a���ƴ'���U�Ѫ��b�A�������'�=Y�_d�x9)�|"n��j;1���ؗ��p����V
u�y�����.��-D}�u�L�(�B7޸�˓��"ĝ"�E�:� ��w�\��p,`D�Җ�x�ڵ�w������aUW�gzxO8��-��b��:�/g���c��(�R��pD�?{s�����c�������d]%�ST`���Ƴ� bE�$�߳j���R��˹����Wk�]^W���`�HX�.1�s䐫�n�z޼H �,Ė���j���%4���0�S;~+�p�k�k8-
Z ����"��s�� �B=���NaI�հ����~MC��X{��l�&�da��1�u�#�G��%{�[-2�����n�۸����buj�[�z����d!Xo�*j�>��(y\�:*�ML����%u�	�dHk`>��-7�7�I4@�R��w@
�+�̫� ������Y�2�z1DP��6W���f�� �=^�"5'�5�D#��|0<��`_���}��0�U����N����^�ہd���{t�d��Y��[3�Y���!)zBkS�(ӕ}T�z\ ��|��;R�SW�j����n�aP�1Ҁ|Ib1�mX�B�5�'��= 3���Oc�d�$�:I\�#'�j���;��Ps$���%�h_��#3����g��Q�Аo��K�ẀV&��� 􋫒���G��FxbyS��j�����$���z��;�<>��ZJ:�j���4{1y�C_m~��{b�]��S���v�R�p]��5=��������nta��Y��� t�V.�~3N�k�m�ݿ�e�h��T�X�Y��J���	B�T��#�|��m��Pq�7+%<�&�_HP6{Ӽ����(�L����h���kO��	J�NгE��"hJS��Et0��˿���8^���ɊREo�n�쵦�������,|�����<M�j'e.��L�]9p���#�,�mc��~N}�B�+�n�-���(�~��0���:�t�%oi�]0<>?����x��Y6��,b3:�Wă�p��<�Z�"���d^�9�r�'��1lE��]$$�^���;�)9�P�� �\�U\ph��3�f��#�c�t�Â&�/p���B�?��>�� ��ёB?�<G��ic���k��|y�~�����:�a��#0���fQCk��8Ʊ95��-�_��wQFS��+��:(�<�a�R��V#��k��;���L���A��&W�'�V�	����홁�Er��&!��A�01�D���������\ͭ�(���(�X�0�Q3���/'T�,U+�쿆9�,� �(�K���.�^�� ���dK���	��g'��:ɟ-�~�©G6�[n�#B��~z�K�ǻ�������ӸE�>p̝C�v�\����0,��ϸj���<�"}�Q��V�cB�T,���K���eLY�3z��H�����ơO�<����{���	kr�P(&�����of���k1��Ņ�|����v2����kq"��R���!��+D����!1��C�S��B��lt[�ͽ������ь_�@9����l.ӂ�'v����0��4����Ef	R�T��\�� �Nh�M����alo�n�)ʑ��i�.��* D���$P�^�[ۂ�v�H��٥�T&��s��;[Md��c�¥>�����0��:���w�Q׆_��� Y%�t�� �FN�(��;�@'�+�,�Û��v����n!���wE�Aǐw�k�r��*�^c̛�c��y)�fQk� ��n֞�I��}��*�J�K��$��?<7<盃�\����	�?�(�߈Eļf�E��17B�hχvk,���Z�v������NURE�t�~��q�.��з�����cIU�YO͑Q�V�Ȟm�s�<�m�i܈�Fs����FL�8)�ǅG����V���Թeȅ����`T.�}�2`�~�qh�L���C�}���o}��QL2�A�AymP@W�opP���;ϧ-�ut�<��ycO��mlD���x�]�E��gi�+����O b��4����wyy���TICt�({c�fC�+�����׫�
~��E����x���u�ʖ�����y�9��^[����[�-®�P/2�����Ő��@/PP��o����v����V��<m�¤2-�]F�����Օ�,z�U� t���aTK��j@��zGړ��q�Jh!s����m?�f�W��1<�H|	>W��8_EN�[�}��X����dSԲ�c��y�:�6�׀���p�^F�����t�W�c�e�����!x���]+�,x+A�չ&i5�Vr^ö���
Ҩ0:E�a߇��~t���ZES#j癬E����n4��o�.k���h���ʰ	�5�zk����?�}o�Vu�Je�}�z�����/��إ_؄s�(�t�r�~h�{��P"�]�����f�H��Zf_�_��x]���H�"|zׄ���lA߰��ۮ���[   �Yb1��<���x�@g S��S�IEz��W����w'��2����3;�������l7���=��A_B؇s @��~����p76A�˳]��ň%#�@'�y��@l�a9бv��y�(�\���cu���b6����Go��ɷF]�H������w�H_����ԙ!�41���}�����U�� ��R��$��	�/h�a��-��r���3g�*ܬ�O�����x ٳ�����5�Ԃ5�z�L__(Eg�߈�K���ɒ�g"�c_\�׉o<�V��L�^z=4_ѧ+��#�<2ﹴ� �_(D�Z�Q���R�x��v���4>t��p��Į�6Q���Ya�h���]i.+(#Im<�JzA��o\�9s��8I^�O8=��+������t$���������AF��ؼ�T�Fܕ��2T[�R������<{h�~��֔w��t&�:[q�w�ҝsi�(y�^&ytnz�'�z��|�e
�1�VJ�W�k��@SY�`c���24�L�I�[L���b��9P��,��R~_	v�m��MK(37#�8������g�:�1e� ա�b��C���}Oe�ɸ�;h�Hr�in�����/���/�"nY���3�v߀2k`�����w���>_��p$��|5U�b�xL���np�
����&	�L���Mi��G���;Cm?y�;��G�� o��;�%B��js�؜��v�`��rF&�S0���U�U�]Hݧޡ���a�=�a*�+a�@2�taԪ�@@dZhS��v�?yn}���i]�+y�Q��Y�W��WTͿ��tݑ4:OP�8U�B���ٴ�j$4�D��$9uU�m���r{S[ty?��s�̚W$3��7u��.ӿE���� RY|�h(Y����ʣ�&gcT�ż��*n�k���R�υ�k�cG	�l�[����&�Gw4��<)�@��O��a�=�v��T��:Dw�q���U�Ta��O|F��?�<F{��$�F�c��V�ުӿ���o�N)�w�L�C:E���7�1-�m_�X�>7!f7Q!·�*�����S|��7�xooKx2����RM}�����[�SHjn�7X'�����|����WI��\L
	�[$F��B3¦!5�<���S��9�J)ܬ��c֠L�	�����
�S� �@�~	ZR�ŞÛ��Q����N4���(e�a�~������lc�h'Ubz�^�~&��#���� ���� �S\�x,z�� �ƥ������(�����Z��F�^�p����ǌ>���1��߰l�m��P�r�M�Q�`�B��)�����C��E19ۅ��\�x&I�����[vt@ʴe1U��9A�W($ ��nY��ĵ?#�_=��L y)��(�	Z�#�`k�-o7���z�i�r�
��p�(�껬�zפ�k?:2��>�tS2Z@K�?=��ia��z]w�c�;�ѕM�N��a��-.����8�i�[�瀢,a�s�E�I����Ȟ'���Xx��骞�<o`�9]�ў#�*"�5�C��R��"���wڑl�i鷑]���2��M~�t#6�Yl�$���T����q�'�	�ji�H:r+����)�x���/�c�Ș)ݑEB�t���侱���)pk�yd�M'�02�F�P�Ȋ����'T�k���߭D%�!��t(��J���@+u�s8���B�n�D�&�"9?òc�Z�8޴,�����> r��MH���,.��m=�������j�Z�p��E"k���b�S��`�U��ᓌk�ʺ�,7S�;#�Ui��Z��/��H������*h��ڝ�� %��@�����������/}�Y��`<nx3+ ��Č\���q�rz=�1dk9[�|&tb\A`B����#�B��l��_o,�[����ʠ=�q�dr���oA�N�|���aR/��P��X��։�ȥ�ˁ5+ֻvϠ��؆�[��ˠ�R�q@��zy�lBI͕lO�ҿ^q�����v +�(��� ͗pDB}�'(:��}�>�f�=_7����ɥ���,���zF�$����c��l eC�e���vӜ��V�#(��GP������jY� �vq{uq�W	AQ�m��V�j��0AIV�����R�g}����2^�V?�VU�H���o�_e[�3=ssZ ��6��d�����u`�2�����/���t%����X�����K.���������ub>��[]Z��J�{sW����ۤ㬂�w��a�Q�*�9:�|�!o��XQV��$di����;��𙳳��J?� #,8�")��3@Vq2:��u&�`���ҡ�މ_>mU�nʛ�PR��1nT�\b�v"7e��dk����D�w�����Y��a
��=S!��;?��Ǹ.A�Ǩ�� F͎�bl��3,���ҙ����u�	b;�Z?���w�?�f
Yi�{�.�
���F��5��*˽/}
�2�@�u��H�b���g=`�%���V�f�6[������UW9�2���C,��M��on��A<kZ:-JP���T;5�B��Q@䵽��v}z���!����j��v��+`z>����t�G�K<ۯ��;�	�:�إ׌V�����#���r��	�폗�٢%8[�0��T>g�1&�R�#.��yls�^��%�u��E��Ej|&o��ڙ��${-4S�3վ��z�hf��/��{K��1��>5�Z�G� x��H Vfٔ�ֆ�$�Pc�&*��R�ة/J��b�:$=:��Y`�n��(��>��r>�� �ć<�ޕ
�q�9A{�����;f:�����M.O�3­	���-BO
�O�(F�/�A�V�\ ���4�����\��� 2D���2>f�������࿄�s�[@�� cB��t�3K�����bN�a?4y����|LT)�TcKA@�BCEJXD!��߂��+&��
s�Ak<�M[nRe���t�r�����u3�+W�l�BOx	�p(Tt[���]�=V�k�`��Ѐ�j�����[m$�$��J��T� 6��*��T�6��B�ᢻn�
޳k��Z�<�s��U?&+ה5sbz�R�;�Te$aq<˰R���^�����X��⯶C�k�i!����
���<�<X��kL�;����!jLFC;V��%р3�Ezs
���iC^��N���V���ȉC�\��N�:�c S7pe����b<�Җ.#�!+M�fAjՙS��5q�o{��	���#��^����5�v��yד�B�i~��ܖ/6�c��x�7`��b�c�G��g��}=	z���9ӫC�_T�;9�)���R̨�x���3�V �yֆg'R���	�7�O�Oy���l�?�ѧ+��@(M㚪l|�ȴB� �Ku�i0� ����u�?5���r����BǷ�M�kD�\&�O����݄���F�X;U�!���ڭ�D��%��1�(ٛc��bI�᳓�yg����e���:F$`��5D?�Qz@�oo�?�0#%o��R��&vJW_)��ls�מ`ƚ�;#���{.Md&�b`���G�dt���٩��0�ā�5��N�ْ$&���!
�_�y9M�+Mz���ԛ^��%[���9P�Wσ�lZ[���#��>K�m�-?`S��=�|$-�`��ew�w
t-o�����4.l��bܲ����ѵ�*(���zP��a\�8l�b_Z�f��g������	���#��I3�:5rŹ(	�%���/�yCt܌t^^|4�bS7=��?��"댏�$�����s�͜Z����x�B�%����8���Eh�	ɡ\���ݟR|��	�{�;�1F����E��X"�kI�Bk^&M;6����Z!|�g������"�E?���|�w
��ϯPy{�y�k�n���������7v4fq���	��.�d���{G�&X R
��ơ5��+��[7�����jЏ��!���Qz��F�!i��'�)љC�ے�ۗX�n3*2��KU5�� �Z'����E��gT�g π��.]����?t~4I�(�6����-(��ȿ�XM\v4��q/D�r$�L�#�Fp�����M�O%�Ml�� g��CF�1�;֐��m^����=���{�D7y+dA�G,
�h���tGSD��tl���4~YqnQY�p󺕳�І
Х�(��	bf�~|��J=�MEjɆp��6�
�U/�h��0[
��O��C����:�%�lQ���	uU��[���	�lȲf�8m�*�����,��u��y)g���9㯷����S�i�i�Y�=�d~��˾r��ژA�*��Sx�Η�E�w!�Vݸ�*���>|��n){�v	j=Y�M���(L
�9�ROx��.���K�;�ϟ�.���_@RxÁ����׷<�ق�$*��8��X�ղY�do�zའ��䕵��/�Gİ�2� 'm�}�᫆X�޵����?��\ϼ1�VN���?0�0�UŪ�A����.�T���R�hk�4�hCI��,n5��J��~�q�虤�<˶���)��y��r�ˑ��s��4A4�{��X�G"O�f��4�4 ºkiؓF�y�i�i���E�~M@�6�_�c�'˿2�uMC�����io��| @�]�Y�V�\Ca?3����Ѵ�v�b���}�U�x��>Yda�9 ���+g)�`�v�xYW�D{����f4k�B��⑫��O��><$FǉM Q�ۉnZYu��^ Zlb�m�[�_���ҩ��uvSX��Wߊ�KA��jӫ�h1�h�}����8���xFB��>}V��Һ߇BϊC��*吝���TM�]�E�{�<� Ȕ�N��JM����L�z�dl!#,�Tpk[�7
�Y�D��Q:�S�w	2-t�cXK���otg�����y��m����Q�i�0�:m�T�k�}ʘ7Ò]`�����Ĳh��>9����K�-��=�)x���v0���ė4�-���-9�A3��5o +�<䕄��z�掶���m+)Ա�%sG6(KG^;(s�����%?���T��>-(]���%�,�Ϛk:����痛=j���@ԬƼ�Չ�d��;*�_#7/T�7əg��m�_����0Rn�>��7_�/��Y�����⥋Fܝ�ۑ.��I��Y���w���]h����|7�=��2����ܕ��:<s(���7�3NȊT��6!\��a0�Ũg�l_HIH)�S��P�K�������h�hw�=Ϯ=���;M�6�J=�o"�|�����#o���c��5�V](��u&���ѿ��U�Q�S�ģv�@͸�]g@��y!\��)�T�C���fi�K�/������G^��&c~�����t޵�*+�|�$>G�'D"����,�W�X�̎i��N�&�ȡ��H�=�Y�+`�1�Q
�z�%E_�^K��աf�qIo����')O�l�S_85�++����W�@3��w��[(�k^6C��-��p��(j�@�3i���l1Fs�Y��+�}��]�H(��L��e�+�Ř���֪�ĩr�I^2%�����b�"��7H��X��Q�㾑�Ȩ�������m�8v��*���Ӷ���Ԉ/>�!qT(ٜ�����D��N�[!�E��8�v��X�m��e�]w_QO�%�0U �x�X�4���AE@<+g)kQ����!��5�B��_�Z��+En�f�Yo�K|D�[I���by�y0O��`������/Eٍ�S� l���h������N�ԅP�  �q�  �󻌎7����aM�{����N�WX��Zb&	I�NG�{k�e�W���,;��>Ǌ���Ю#9��[r�T�ՀJƆq��X(��aɇc�_��U������
�=6�����,�SLR�0��u�֗^����jI�0�b�Z��ٛҠ6!GH���\,T��|���=�9�3̴ʕ�I'��N�@��� �����*438���bE3���:xҠ>�������b�4�ц�p��*�@Jp1I����_�Ooǀ�x���`���'4~�pgΉ�$ozF�����o7�);��Yȉ�^�Ε5T/��>���R�\�;=h�kO9%O�S���X�|}�?Zq�}K���(K}��lD8Q��5��V�N�޾���W��'�R1���J����~ğ��4k�4?5Xt�Fu�s�i[n�|�Z�	��~n�|���2Be���ϛ�T.�����^
6�a�~�T��a3���8�0~���%�&��Ya�bc|?���6{!�"~ �&�u�i�z���C�Z���9�;�u��y��R�ZD F�s�.Иp��s9%����E	��;H���-B<f�[(�}��K�f6���}��	̟���I�R�*8a�+yH�����{ �����I�Tlx���YDg���PH���,��^W�o��W*�xe-Ա9j��O=89�����~WA8�_�!9b ��i�_p_T���
NE��b�6�j�W��2�k5ۯ4�,xP�'n��P^7���}��~���3R�	��S;yE�8{Cc!72�j��cs�����*XUf� �g�5��Qqp�U�)��(X�p:O�T�XLn6���;�}��-�p!�?��BEg��_7�O�U1ѐ�1�b��C��a��<���z�L�����f��]���Kiۖ���e�|�u���!��2b��D���~�ˈ����%���^l7��_P�o��)K�׃����O��b�Uk1ZFڲ�������1gô��]�e�}��]dgF�
׍Xv����j�J4�F4GO��<�8r�p��[Gn*�'�1C�� �f���R�����aJl����.r��*2�Q�]%�Zo�&�$D �c���������jjl�<L�;��v`7�?8i�B��>Ҹ8u���C�\ON>Z�K����k{kd�$?��~����gK(1g�X4��W_�����o�j}��z-a�$���?��;N�'��Z2R�{���a�PwT����q�o��Δ��J�c��Lu�Y@����Uf8޺(s��úG�~�#!�͟~nS�v��b�2���2�6��n >	��������.��ʚP����~��Җ�FR�p�F���ך�[R����j`��� ��e�c����`�,��O�µ��l
n��>_K��}�ӸM��v�&ԝC�����`NZe��'	W���I�?X�_ ��+��6�qL�d�Χ+�k�"u�4��ut��"Հ/��o=���eꨯZ�GX�>�������3���4���P��h:��Z�z�m
�+A�~A�O����m��mg�9!�~�M�$���s��y��{ˢ�!n*oR����-���THA�ߙ�VCnOU������r� -u���u ,f�rx����H�J>����L����u��2G��'�2iq�=�^���>��,2Q���F��)�d�0�D���Ǉbٖ��;�,ɵǫ�����`E!?0�N	I4���(_Q�u{B�}�bݢwAT���(,��y�7�w�+�Fs
��)'2�;�1��_4��Բzx�a�Ր��^�F,�.���ZW���y�E�wy���y�צ��("|{t�Ek4fm��84��*���+S���C��8��J�5(���]��R�D��A������6j�-4k��Q�l4x*�l`Y�d�1�Q]%����J�Ԃnml{݈�G��'xݪ���b��_?o
oģ�Vٳ��̳7u�>�@�5���:��j�,cZ��#Dj��q�'�����\@>�\,�7����ئ��(>�9"�}EB<�Nq�B��I�Z�mym�foB�0y�9(o��2��w�8O���y�����z��q�����@ >�wK��h7T���$7������A�:�צ���9�i�g�ܕ��P�s!i�17
�c��Y�O�1z���R�|�Wp3��+-��m�Zޣ֛�{~�4je���9�yE���z�,d��U�k�C�O�GZG:@�b�^k���_�m�ƜZ����ͱ�+>�1�	�)M�+"��]vI��K�>�Q+����l�	��({��ח�Sa#'"��߁E��c���7�q��-��k-�hlՄssS
����wK���t��e�|�HE��%�A��)�j�w����E�Wu�v�XZM���,����`�E��Y=6bC���	��_F_�$��FL0�K1I���#p�:�:�M8�W�7�1�.������&|�LX��Ύ�1�6�S��uҴm0���x��B��t���
�j�	�ɛo$J(�j�����m��4č���T��ĸ���W��4��M{4/$�?\�����V^���~����fmz�Nc��|�6q���g�վQ�@FxD)(�����z~�R�>[�)e��%�
qL"��)��� t}+S��BX`1�l������b�������͹�Y�z�!��f4{O�%��ޮ��2j�[6_2���Y�6����j�*$#�K���,�C՗q_���"��m�0=3���n,V�R_I�3�� �N����Y�:���Й���:�+(3/��IZ��F�E`�lkZ���3�j��(��ĳ{�M��1NǾk�h�.&��y%18�R	��	qk%q��J�?��h�{�$I%�f�\���{�4{����\��P߀u��!�]�!�%�q��Mg�"�+d��DT�pR�0�����^�Yd����R���F��j&/������f��m��DP�$�-�HcNW�`+Jc��O�,7�!k�{�Y]�Ys�N�m:q��4�\*2J1���-�� �R��&3ƚ�.d�u,�QCy��Q�w>JY�QhO�cXr����i	�
��6SQ�x��X`�}���A|lA㝡��9��6B�
�a\a:-�I��
�Õ/Y��C	,��l��d䡳�T�E���I�U��b��9@��m���0���(S�-s#��F�6�i�b4��w�Z�EA�]�0�/���e��Ϲ� ɧCh��ek�u[�\���7�UR�â�XZ/6�L�Wi�0��4�
��\�ٵ�����e�.�Ē3�� =��W�+35ĕ,�;���ۗ��ȷ��fQ���E^��;����t ze�z�U����P�$s��R�nw�Ñ�[}���QjB@K��=C���4*��~�4�c���r�X��x�OYmٺuv%�����}ʌ��UE5= ��ot��1Y�I���9gB��X�. �Z��bX%���݁w���3���_d��n' p_`�7��I�0��6�'�a�C�mȰ�U
08�K��iH�mo`��FŴ�K�n$:t5�)?��zɒ�]O�e�S�P1n�<�Nr��-��M75�D7p����:?��j�x<���1Bz�5��^�}_X�ѐ4�8�خv�9 �Nr�"^Rf"�!%�`�9��S�u�oL������Y��'��u�C�@�@�{ �s�3�h���;9�cC�s�S���ηE��[ĭa�GE�����|̺RJR���dw���A����+�؝q��C\�CO{��3=-�7�ɏ�v3���l��WNG�O�C��2�	�=���,�s6(=�mAjbg'�>��~�ɷO���1��?|�_�|Bs�P}���1x�Ī&��$x_j�5o��l0������	�\�G��f���gh�#"�vh�C8��.�+W_P�<A�h�T��46��o+6�!Ü�5��� k'Tᆁ) ��jLJ@��v\2�FCwݐ�_�GϓR|��%�Q�Z�%�5&0o�`�RM�g��s?��S�&<���f�˰���3����*wv@���ԩ,�[��in5�*�B>5��V@��5��3L��k[�YΊ�p2C��ڀgQC���!�R�]�7��)ܿ�;h�H/66�L����f���R�.^KyPԸ���
2�K���!$�G)B�j���=ߟQÂ�UdX�h���e��T��1����4j\�]��pDB��i�M<g�k�����R�S?��(<ۮ�Wחh����v�g@.��Z��G�H��&{-;9cL�+�	@O8+�U���r0��mS���[�dbWG@�4?��*O�(�W|-6��pJ����	�ЕN�u�/2����F-�%s��{����xz�z��,�"�N��
ӂ½�g�՚K�D~y]՟w�`��TNRQޚڠ6Ǩ|��oi��i2t���	��e�$�(���� X�q�$��5n�lU�PK�R�F�'a���	|M��RbRլE�Hm;� ȯ����e3��-˧�Ny�R�ݸO��G"�w�)Z���
p�P/c\� z�Ž�7�C)ז^��`�Q:~;��5.ڮ��f;v��#�F�}޷5-"��C3��fb��,n� �60���X���Ncf��w�9�m�����6��-u���7w�x�����b��L^7�Hv&h���b�Ʃ^�X�n���ih����X. ė=�SC��4�_x��<㔠�V�hJ�(�]@�o����Qu}���.�� i����� Jw��?v���U>�f��%�R=��	��V�;Hxn(;���HD� �s��ut��Syң����D���<h�,]^��j$ঠl��f�_�V1��7 ��SG{V���
0���g����|" �
�	�pm��ǈz�,��Jv�ZY]?:x���؛�fgJe1he� �VA��ʪ�+�,Fz�wI�`���)�R��l�G� ,<UE�H0����~�t_��3H�W������Q&����S���C�=�t��ɡ�W��A��S�GH������+��IS(30_���6C;��n�'�,C�O�>��<hʌ������7�"[g���yH���8�S��&6n˚�;�Ռ��bC�a�Bei�s~�d��0=����)*���PB�lo�Ȍ��G�O��C��5�.��D�������y�[`����rv*�oٓ��t\!�I5z�L�O�U��P�aXUex|i���{/3+��\�4V;:c�F��þ�p,�~vS��B��ANUu~�2�
�w��E��9��I�Dz�U3�P��P0�ڛ!g8Q�/���e$M�)�Jף��_[�8�����-�9 +�'�_eQ}.�S����^@_�8�����D�a��/�Ĝ4�5�H�o!8a/h�wŵaN@���0�󗛕�;n�/����e�}h6 `L�)_p��AEG��!��`r0~�Z
ҋ��-cL���9��������
Lsx�8&%����53��E�duz]�a���`f���*��x��p��q�Z�=��x����A�ai�7�*_�㠔(%������-d���"?�2�́k�˩\r���h�\j�v|���LeQ�"�����O��Tr��$d�n��$���5	�m�o�	�x\�m.HQ���Fgk���K�~��p�v��.�ZN�|�޳�cU�����$6�o��֋�z�n���B�bj`m�@��5�u��Ó�y&s���UH6�vv����Œw5�"g�����ն���쨎p�O�'�%�����l�s����y}�r����&�����d:�Ǽ�m�Z��ù-�ni(]�˃eo�q§�D)3ٚiP���0L%|HxM��06�-�Ȑ�l(P{�啣:7l���R�]�Q�~`<,_����9�k�5ט�8	���j�=_�!��`��*��O�R�T��^�	i���7{�$M7������>ݫ0F�_�/E�ˍ`lz.L�m���b�a^0��Bs����Z��_���gR�~t"�E��&�����z��^hr�a�мA���r�ja�%�4��|bq��0�t�Ѳ�L�hr����:�z��mB��"�m��3�4�����k蒂�b�;Q+	�hU�S�X�}��� ���D�0��!%�Թ���=sM{%����Gw�� Q��~{v��d4:���kW�w<��1~��{Q��%�H���´�Y�֓�H:���-%���k.�,a�����2�~6l��w�N�@6�գ�M���z Y�ӿ����8{[']�'�)(m�O4Y�z��������M�v܃t����̳�Y4/��(�{qs#14DL�gJP��Æ/��Sd��MmG��V��'��F5g��+
��~��#��I�w4�#М�:!$��B��Jyy�$�>ʃ��ڇ����p[��W����J$�1{㕭�5I�3��sÊ�.�Y��O�Dh�����0����l���^79c��\�ň��3�����FtG@��Ke���?�'HV��>�K�6�ǵ��9��E�I�Z��F*H=r���%&���1�����ܻn�+z�R=�9�y��'��[�2���,B$�=��AN(�m<t�E��O��0Jۈ�F�3~�*�]}�t¹�hǮ��c��R�&/Z�#�O}]�Ll��ˡ�V���I	P�(z^ۧ�=�4�tX�	�t�˅<��n�X	g5�#�`s灭+U��XU��So���[�#h�*O��/gz�fY�+- ���G1�J]�H?(ۜ��~2AZ�7��ӌo�i�N�C�L�Bj�"D0�Q)�r���R
5��ޱ�Wn���������>H�%㷺�uU�W<*C��g����4Ԇ��5FVN�~S��� �dJ
��zb ]m^��ZC,lE��*�6�(>��A�Y������>��h���pb��������g+%�d�� 򯰇N�V���ѿ�*�~C�$ߩ6a��g1���Y�]�D����
$1���*~���eR�8�����XE"T7ɫ�c{��/�C�Ϳ�6�@aZ� �C)M����	�MB"88�r���ҩ�o���N�@����]XC�������m;��%z�DOٹ�>��"+
��v�9��eE��e������]A^�F����,�\G�)��Zi�ڡd-�Cx���ǃT�k�ta:E~[�ƪ;���J�XT�:O��L�}=�'�V=1*��M��]zddc�5��qA�"��:O�o͘�_�|w�ŘT~D,
KlcSj� �p1�|�)�72ڪ�9rE���<���3�l>r����S�������u�|;H昶c�U$���:��΍H<��ۦP":�?�A�J�ܡ�y���G�H���4�Y��2��,"m���g�ހ��n%<}�N�G��*�Ȱ�&���@k�[���W�l��}/�*k�K^+�;�I���'��Ch��KkE�������.�(��V�@���ƶ��ElcO.]5/�z�Pn���� ���.���]�̠)i��?�k������K-����u�xe��o���ur=6�>�'��ئ�~Z�q��T3��'��1�T~��p�㠥���/����O�,��s��F*ˌ����3a��62��؛����-�nP��Fi�	G�=s�R�Ʋ�4�b��w��6���Q5� ���;"���=ˀ@�qET5���a�v�x�m�!0��"�!�<�M](���!0wY�H�0Ao�f4��p��W�$��*o���o���Z8O��J�v��
0M;��x�n]J(�L�(����7�dؠ9Dr��Y�:����fx��n�@'���y,�%�5���6H>dR΄�����f����H���W[��_Ƿο��sAy�ʈ`0$�_��'4�(��F�	�6h��9�ܻ�ھd�\��<�b�>�ZK5;0���-<�3Vt��Z�`#Msk��:�
�E���$9<B1bJ�s���UD�-{0�I��X�u��x��?U^B]� Y���^��0�D�ҠZ��?��u���q�G��!d�7����O�o��n4�Q�@�lL%����ߖ��n�-�%އ���n���������ؿ�٤�)]ބ ��A	x�ߡ.��s.�X���`[�{p�[��=�ߤ�C��RD���Ib��62������`�����z�I�9o�iь���)Cc$�2��va+� b����qvH�N�k��y�\�L�ɸ��lIvF+r��d3l&\�1G�N�C�|�|�N�_j%�q�oM���TD
� @d�Y��Y`��D�Lu���t���S����>53��!&�y �6���{�U]�ڹ)Q��Eg�������g�s�(AQ�c94�T-�W�{oM�ޔ����'����`
����qǰɩ�~(��/�@<(
�$>��I\\u������!d�,���0��P�����Y,��\KG��R�U�VZ�Ż[��пm���X�L0�XI$r��m���»,
"2m��J��R�W���{�9����9��S���$��1�Q�8?�����l��yt�:.��w[bQ��L0σ�)qw
�U��\�Ms-��ܠU.��Tԙ%��6�fϑr5�Aع�!�*V��]9h�6?,�M���]W�u(���q|`��`Dč��ak�Z�k�H��챟O$�x�i,Jِ�t�E|�;nP~1���c�P�t�Z�#�&CÕ
�g���-L�?���k�L̩�Up�sз��jx�9='j�]450��/�h�߂�(V���S�2E?F�l拺V�8)��Y��n��k�f� �4gsv1 ]Wڐ�b��,����z���sÎ�v�DH���D�'\]�K��V���2K�~�9o�F���Da����l�9�&>Y�aH�.�
���3�����l�
q`Jl6�aZ+�)�;�F#4F�|����[�x0�a �\�d�r���"Ȫ�~��-d�x�Y�����rK���U����-�c�p����������`����� ���R~��Nv��r5ֹ�o%��{�7o���\פ�{��m�I)ה��m/�tl���_*�$�v�Ed`�E^����E�O�t,!p2C�>��p
^��<dR���*x��9�h}��viP�Pa:��B�s�O��&�Ys���ȍ�Z[�67,�J	9�
Gx}���^��랜0���}3�v/��O��J#Ǭ0c���ˤ)�C �?	���`9��ݾ�m���5�$V��Y�r��e��jo\�3�I	���+���5��6�(�?��r���f>.2�臣�V�CX������𐌙�U�XK�D9�R~��)�L&ϕ���ھwPw��jTA�!7��W�u�/�z��Ngj��N�/� �6��k=����~��e�^��|�p�"�D�ԜȄ��kN��z�A���},v'W���9&�6��0�ng5.T�[\�_{0��=3�Z��-_8 m�
>t�M�?�i����xA������
w��E�j \�?��"��(,4=�ųnz���+*�<"�dc`Z�"�蛑�.9\]5@�`Q=� �&f&*;���+�Hv��>�]��U�j�]U��Ei�#�^"`C���L���o�a�	N�����������ɀ݈V**H��q��\�m����k� |tIS���̯���<=ʂ��{�c�Y�x��+���f8	�]Hl�?����D^�L�;�eU!m�@���T�T��~к� �����025��93�8ǝO�H��n��vI��+ZF@(T�%{�ʲ%�[�j�~D]�0���:;(.�� 9|�A8�ĕ(F%<J��ҟ��K�*٠*��v��!�**	��c�G�3�/��_z�(�uƏ3���~!/�j}�'�յ4!�ў�/��ZC΋�=~/�!^l��/� F����
��C[��y��]^So9I4~�ᵝ��r��'gT8YHI<O.J���%M�pC��X�h)�|x�,�P��� ּ8Vrx4�t�"w	{���l�폚!���w~�B0�HXh7ܑ��y%�&ս�l���i9�-z઄��X�k��b2p�U�]���/�d<�9�8��{�B?��)o�c''�����S�o��u&���=��*ok=��l؇�Q��{e�����J|����8��)�}a��q/[�h���������z}���H煛���jz�-��r���[ߦ��ߡh�BlU�:>Yd�$Ic�ɐU�؆����R���mq(b���䝅깈@��Zْ��,q�9�5 v�[T�6�T�΄�^0���m��d�
̨�P�P�	O�ɞSQ�e�� Ց���u�J�Ͱ��{�BG7�Ⱥ�w�yx�H�һ���%N���S���e�x�����A@�n
<�A-�q}*A��4y�b�TLп�*��D�ZE`�ftP����8 ���yP?�&�la;�tҎx�L�xA���ޥp�"ּ�o)�R�ڦ(��pё����C���V�^�>�@|��d��톦���*>�X7��DvL�����r�r�k^H�N&�#.�Bo��
�u��k�T�o��o��Gx�H���lr]�d�9<l���\��)v��0��	�P?4U����d���H�D;��f��ڨ=i�y믑|�{9�Aܵ���䒷�K�ث��No6��A<�����\;E&���c��T��ۣU�o=�ւ�|'&���>lq�a�g�r��ޘ~�}Kx�-�DD(��v,q�l����v�\�@Y��؀��8�>ۚ�g�m�8������_h���-�\�ue(
eQf.3����,���h���5��*R�ظ6�S�%��Ȗ�8�!��S�w3[]�r_�����RC�)Jtj���i3�1�+N<nJ���)����>�+�(�3)p���J��^N�����TGo���[��\���͇'��bҐ�^���@9�d��)�p����)��`���)N�8���J:�~�\Z�69�L �*��z�a�	��W:co��Tod��3��gk�t��8I�@�����Hg л�^��X=28�_���Y����.��
ˈ~������cwP�g���w'θ�ͷCkf?m%`<ε8~��WF�^F�[7v��Ѕ��euQ�X��j>߹���?S��6��Md�F�=?��Ay���J���c&�R]��X�����3יE9���R����#I��� |��/G~4h��`co�ĬL���-��������
@��</�B�O͙�$ό����I���B��3������G�:F����B�����ۣ��s8���Ē.>����,:K�����o-t��zF(G,��	<���t5� n2�[)�["� H2��M���6@���Xj���n1D���m�	�_ѐ��m��Z� ��@`9���w�)\�ܻ$eP��؀W�����g�Ws�DM�v��-�̘�,�Ng��!��N�'fyW���K��äa�E��ms72�wY�����i�.�j��$���;l^ݾ[�������P�������C���8��߲S,�>��w3����R�J�^��^�4fBil�>4�3.aN�B�AB_N"�[��.�	�-��13+Pup߃	�����ִ�w��F����\����5��/�D<i�(��v����p�UsN�g��ka84�i:.��eLD���{�=	��u���qѓw�AF��;		x=vy����_�J���L�w2��n�T֣6�']�z�WJ�MJ�͙���z�B���ކ|��WQ`���(�QsQ/P ;v�HR.X�*nA��d���nR]ijf=f<�v��E3�Vؐ����BE�R�.�L��K=�)Ш��Gd���gD�S���!�4�|���00��Ĉ�o$�F�� �G{"a�.%��<a�ǎNp*�2��� �s�Q������Vl��vhL�y7��İU�B��E��������^�s��}��O�Bo��d�-f& ��$4i�m!R��3�D�oUO��rMr\Y����� u7B�������BL�R�)��`�isr"'��t5�9�PF?o�������"m\���"�: G��h�����ڪ��ST�!�\��gJrnZ�Oo�A�p�%�əI�Ng�+V�6�\��ݠs�'�,>bV���>�Eg��x��n�A���#1��Cj#h�
��"vj���ٸ���X�B�/��!Y�v[[2묶���lr}���-�>;���+@���ꏌ�t&��A�-u��)c`�ٲ��7ḁ&ٳ�k�*2#t���p��B�������WJXX5��+}q�7`�%�{��ثƇ�v5m�L,�3���1',�~��q���:*�TGؿ,f�X!����5<[��|JRՇ}=v���}ý��w�3C:��1H��AZC�}h}����kn�4}��+�u�w0�hPg8&����gB�"қ-[%aP����?ƒ&q�{�>���	��!c+���6@N����4A��7��n��;���+��7h�S�碸{N�d��i�-�F�t��9�'��_1x�1UH^VLS%����=�{ѯ���BQ҈#�`�%���n����Y �O��8�Sn�u-V��19:�pr[�h{���
,��eB?���Rđ��Z?�������e��rʂ@���ߒ<v���>��fM�D���Wi��&^6j˪�O�)<�:6�)��B2�l��bS�Oi_�S�F�
i.�_ a��@���-)�ɴl��;!��p۲d�'R	�4H;��a�t��q�X�}�%���"y�nPk#�r�����$�$��w.�qliI��ː4��)dA}L�����j����+����p`��\F�?�]տ��,5[�-0�x�̥�b��}2;=�E��?�<��� �9��S�����v�B�l����t���e7Xݭ������;�؅�uL�~�KS*�\:�ωGN!�@!�Z�G����}\�G2�R�?�pT��)��Hp	�^`}�gB�V�1�]_��oj؃{�s�]¢�%���?�[nQ�C�E^ܔ5�OEE&Cbv�t�9���;�n������<���_b�m�6�<;��K_�"�*6�8d�&�o����q�+�Mm�2�A[jw�����AqE��>�C���crC��e2lhB�,���2%I.���T�%I� ��#%K�{�ڨb��\��Z�k�)��eCO|�'��04�㠸�V?j�����it!�͠���z�?8Y�$�C.��z��[��>���U��h���o�fc��F��T�����:�H�M��/b����X#|~B��R! �u�lc�N�N�n����Mz�&�	�wy�}�����eG��U�0�����~w�E�6�_��z�w�`ꝼ*� |�y��s4�N���3�!c2��V�:������ޮ��N�2�_�\����,a�Q��:b+�x�5�ȏ���E�<�c�fwG�~�F�r2S��[�oWݿB��Ѣ��"fK�d��&4��y�p�*O�ɛH6�ݩ ؐ�1�?WA��1�ۇ�:v��ci,Q[8T�U�u�#CfVK2\T����mL(#��u��B#�;K���Z�� �%o�Rbf,+Z�3��t䝝��L�u|�4Y7<+�̚�_�.a�pL-���Qx��悙(�������$����BK�L$YX�ϰ�ſz�)ÔO
?�������B������(Rn���90�����(O�4�P�x�`�����/�iu���c/��x�:Գ*-��]l(Da�R���a�i)�;�=��v]��f/�{)m ��>��o@VgK��Za̬C���	���Gf��Ł{,T[�&�o}٬'�cEhޗ&��XU^�A��%�|g��dm,-�N>�qǎv��=*�Xn�
TG�$�p�OK!��s��d#��Z�r;(��B�Ik�L ��G*e��21uOQ�������=����P�Ê. BB��f��/�&ͽ���m�ZU~��0�j�K�EH�����S�8Q���k[{�4�T������=�qf��lB9vC_dѰ��-���X�����<�9u�����YVxo'��n_�i&]�z���*���L�p��f�h?J_an�2q�qaW>�g˖�QK����;���lb-+���q@Ơ�-� �H�@t��!p���!�:�*�����K}7h`}�w�����[��K��s�/�ɲ������pn���
G˨\�K��������^��Vu�f½�e��eY�
��O�(3˰5Y s̖θ�#	���e��"A%�=�Q2E<�m:���>]-��t;�I�?̕Z3sH�!�v�r�d���^�V���e�.�
�	)�Y��JG�?�+ģ�DO�������݄pۢJi�ɳK��UgH\
���;0/Ps��*Q����W����_�4�mB��y�i�����/Ӻl��/*�_<��H��-���)"=�4� %M|�e��ګ2Fo7�p?F���ĵ��\�#�ܗ����Blv]2��ĺ��#Y��`z+X���zI�aiW�?)ܵ0�n��Y�a)�n��SZpP����[S��Q���Hv�n� vU���q�!m���I/�4 ����5�x�q��SY	G	+�["�T�� o���^H��i�6,�D#��yfc>oɗ������-�gL�!N�T��45x�L$/�*` ��e߂Z��#�	�]K��I$6甮������������z������;4���oi�m������hD:1�8��;���v�TW'!w�q�DJcR���ʎ��/����E��5����SA~���̜���O�i�����`��d�k�OQ$�Kٜ�xe؆��[5�'�J�o���|++V���߇ꆈn}
�.h�l���#����K�.�R�^r� � �s�n��k����bo���Ì8�%lM�F�N��N�j��K�
/N��śx5�a� QEd�rV�~����\w`J�Dt`�"~=�ۆ�d���l�����B6X�͸��9�5�St0Ңz�Q�FM��Q7���Xs�6h��� �����5�t+�����I�� �*E\<�!���N���a��6I����E�Z_�8{���=�r����x�5�n(;��*#�Z�sK5H���Q#@���&1�ѝwB���ȿI"�D|5
,���s���O4�OE�p�yGexF��H��)=lQ�Zˁ�n۞Ν~���G�U����Z�HU�����u"yH���(W�1�Rk�2d1�����:,\H/%W�?��qj�i�6E�ApŃ^p���sAHg�E%�UL�6�*��~F���b6���_/��h����C���G��U�!�=���!�V6^f�3+U�W}�p��B�����L��%I������"��#��¡��x�?!�%�UƟ��u�g��_ZV}�$,�����AV�7#��\�g�.�D�f�
I�	�wX���Z<¢0��´Q<@��L�U�J��4�W��=����u�lW�"�4�̸��Zm.rFىs�2�X�����3_1�wb�n�Y��Nm(�i5��xL?VR2l�H�z9�#��C�5��>�sLDb1��,�vZ�uyaj!�@�o�rA�9f:��$M%<�SYf^sΉ�E<�| ao�?r,-Eʄӗ�C
 (���k\�p�gI�^�i%)Y(%iLy�DehM�X��������������-̶��ٕ��M20:��Ӑau�3����<��b�^6Q1�1Ҏ]��0$|��'���Ӳ���nS��r��^d��@7�~�6�%��f~m�α�Qh�UyF�K�F&�h��?(ݕ�)�K�E�u)��>�o)�O����[�i�<�9��\�����������Y�z9���x~?��B�Xt�����MM�Ԗ|�V15���T���d�5F���: �o�����������Rhbد�,EֻDkV)��be+kt	�P��6=��*&�4�v1��}������� �[̑b��.x������/)mG��V�|Ð���s�;���U �s��Pw�ZXs�Z� �	��RH�奀�%�NͶ>w�򌲽gwÒ@�Q]�u�i������J���N�����p�����K��*���e�<�)p��O�����J�v�{��g�	�0h�^�Y.KbɰX�{�G�c�I8�.��Vh�\�0�w?K�<��C[c XϙA�Mٮ��0��L@�Si�|/My���o=�p�5O�_�=E�+����޿�+H�&ȧ?Alf&�1��)bz�����7�dN��Ν+���?�olG�v%l�Eo�ݍət���UN�2[�p3l�U�C���OZ����nM� �<��[�7j�-�t8���V��%T�\��w��,B�"�/�N�u��|�yKB�4�.j��X' ��E� d�6��Oz�[V�o�|]!f��Iu�P�(�-޴sɟ!M3�����[\��J����=s��G�U�����$_~�Ͽ-�t<�a�v�eDbb������λ�D	.<Ar7��4EҬ/{��[��q�U0�[J�ED<�%w�oB�˄a�E�R3&l�|������O�@q CN�h;�*9S�f��-�S�����n��YG�aGZ�-Z;�4������R�"���Ή�(���(���~��`�<����Ҫ!�)��❉^Y��F��Z���K�Um�k���_
-{�+c�Yh��KdK��B~�Q�?�By�T��D�Q���+�'�Q`�/V�"G9(?~��B��H�o9G�:�:�&>�C�x��ڜ�c�s��*sx5,r���+�Pæ�Q9 Kx������:��d�\/i�s�@Y8����O��o��#'~�5��3z���ؾU��Eh�i���wXowƧ�L�T/R��\�eE,����_#��pJ)�ңk��^rmd���G/��	̡���h��ǥ0�ց��>����h*T�]%���/�;�Μk�<�V�6L���o6�-b*[�����U�����@?S�
��Kͻi*4T�f�3�:G�U��q3���zԧ�
ZJ����&�
���ċ����%�lr6ds����0f���D�sx����-���\Q��.Iʩ�Pi�z�Se��5����za�݊��ŕG���_e�������C�U��4-EL=O.�D���HK�2E�9-��f�8��J�d�rH02�_ ����Dh��h�b��^^CA�v6��#���N~l�$��.zCR��'�w�[�:�d����?�М7����r/@\{vuF W�gs���VJ#P(\�\�0o^���ė�m�g�C�bSvXo��v�-��יH���Lqh7?J�_69��x�/R�r���O�,;$���޾��7�c�L*=<��ȁ3c��z ��;z��99��rI��[��z����:j�k%��M��Gf/����hW�(���>P ��$��h�m��]y��qd>��W��F�ӹ3��Ԗ��O��X�v��#J����T�$~׆�!V '3�� ?ujo�Bx��N���N;�,��xW�x��
��T��WI�s|���Ytu�OI���w�[H�n~_�1�x���!X5FK5�M@C�S�ĪE))!��l���wi�!^��^�r����(I	"�:�T�=�{*�:��ܒ��m��A�k�.�� s�o�*��`�h��af��^�mgrb�nS�np.®�K�e\���˩)T��� ���C�f|��N������h�.�oa��}����\���KSD=XJ�u�����ј�NX�6; $!�Ά���޵0b�`���_U�(�wnv���|����76Ȓ�0I	*����Rjdw�sy�G��*�1�)�d��~�E�ϩo'l)��#��N��6���x�P��� 4,N$&��|���N��,�Bc�pY�@ϭ����0Ք��e�v��rk�ûE�yz���"�l{`�P%�==%$���8���gL�p�n|�h�&Fc��_�,�~������mB�)?��?��0�ͳ���%S�V�ًGy�u��Y�rCE	uK����\�Z'�?�Y�zϔ.:�,m�y����F�v������&	�]B�[�<	p��v�O0nYN��do�{ir�4�i3]\���qD<oG���~��h@͹��[���c� �=aJQ � Y���ު�K�g'�^��m��ɳ��V#��EV�fy a���zS�ߙFa�+"E� Ƴk*;�GC��UD�`q�"��͵��y	�V��^O���F�tc��yg�D���H�76�RGq0�ͳ	 B]�E�1a���-�`n���ū��;y�*nC_^'P� �N�3�,��K�GG�2`��\��8c4ZB�N	d/SK���-�	Bӆ��|�`�𦕡Jyn��t����kT�6��mz+LdQ�*�ݎ���c[�ۂ2Ȯz����d�dm�b!DGv���b�7?T��6�h]�5B$!��C�'���pi��=�"�6������E�4�i݉�t�`�A���dL3��k=��#��%#�`�j�����6�c��|m��Ԗ�3�pi��{8���aTVO�H6�<5\���!c� �/�4��U�s@$����a�Sl�)<r/�ǘÒ/6<V�8D[)g��
"luQ�&�ii bO/�u4�%�jJ���m�f[��Ä���þDZ�Ӊ9����6>�A0�R5Ύc� z�n�4׼4�*P�HŐ�0U�xdB��b���8ᕙ�Y��o��?hk�\$H��PB�H�|�?�?{�:R5ix��,���B� ��
��<��Sg�1v�1��B�{������T���V��f7di���N�乺�h��X�
�g�����!������Oq~NfD#,������1��,D��ӆ ��X%�!�_���~�(�z$�	����h_���ҙ�Ͼ��H�|���0������|wX�ކ�sѦÏ�4:&�����z`����ʣ�mt{����A�ɠÔ�A�2����2{_��`#N�+.��
����&����3�����1U���y�\�>��y��q�!FsB�-��,��W��ռ�5�6l{��Qق�t䁖[����[QFKĤ1��8I����Ĵ/r3 nmiv7�<L�����(xt.��Mv�6���f�g6�
1�O��x :���+*��
G���L�xX4�N��<�Q���Cp���l��
o�����3����g��Zc�}!WjsY���V��t+�8Ɵª�~�	8��7L�w�5��	�z�ז���s^�45�D�Ӧ�
?l�I�)X���)2�ъ��t�vtYZ���f�[_�2�������D�/����X&X4�/p*���
ƽ�
]��)���
�lJ��x]Ī')��CA���˄����\谟ۛ����_į�Vтj�v�P~>�U�9��b��:=ôH����{�ĲM�3�~/]{���!���:[����M��\��\_Aa�RB�8)��)�YRۺ ���5��ʢJ��Z�e�O�3%g�6��#���:?����������kP5�c�R�������!L��yC��o�� �C����Ū�7݋'8��ԠU�[�[N������6���e�Q&w XH|>J�h�CiB
�+` �Ω҂��/���{q���j"�7�
 _S�DG�=�
zX��c7Ϙ�?�=L��F���D������X�a�Y���Sp��&�iI��f_), e��4XMd ������@��A'�9`	�]0^�r��q�b�k��0��XЧG��־�d����j��Z�
�<��C�lLXJ��b-+�$���4uQ@E�i�ɫ��n۬(�@t�hoy��ǯpr�.�A��݁��/,�B����c�t!�7d[(����/^say����D<�5�C��e7jL\����{�#R,���<C�ځ�^�QN�ri��̗/�@ny�v�@ߕ6´�r wA����=�P�h���0��.�9Ʊ���(���^^�&lH� ���N�o����2��HAC
1������qwi�!?�@8�U+��*;7DwF�5+X�ڱ��l�q��D֏�f/o���.��U ֫�n�H�^�7�+��)�'�P'_���9[�3ƕ�y
d'���_K�V��\	��]���~����w�������;�O�L���`������3v����l��*���.<Jj���N�6�"���&���[������q_ ?�#T��	Yo���@z�
�{�h~�"kːDC:�����!��bb�rL�F���'����̙�X��;���0���p��M `���<�r	#�?Fޭ�S\_'v�R��E�ײ�g���l$���%��A}�4KWZ�(U`ם(�su׬tɷX8\M������l�R�3���kFI���/��0�`Es�)�q��&����t�[z!�����ϴ�#�P���zjr��Dd�@�H�ߝ1S�^��8r�t����Y6��/��e��Tw�3"N�|�3*؛!`�6�ē�3�{��x|�jç���.^t�k���$4@���7��i���y��	��s����M&�R���P�)�V�N�7����� 5Kc��7)iV�B��Z]=��x/wg�=�DK����c��x�$h�\Myl>�.cV?z�����&�9i�0a�b�	Zf�A'��*�('�S1*A���I�W~
x���q8�8��(��aH�2�c�DQ��H�L?±��-��*|zÑ�]h����,i+��Bu>�a��F���K�,xc���Rq�'����O��X` ���3��&�fۨ��ؖ��
6�l(��N�~��Tݜ�}>�
*��ڃ��ZƸ�(ݣ�^!�}eqO���@��7A�&�[���[�˽��1���dZz��̐��~���=�̌Iw�e�D�J�\e�-3WP��+ ���^ ��z�s�,#���q��W�ƉC:��8��_ԧ� ��efB�m6�tl��D�Y����h��2D$����|zEףG�!�����:Љb�0Ff«J�b��Л:c�0�����DN�`���	7d��\nҋ����:R;���}4����Yw��@'"O0܅fX�X|0ɘ��1�'�c���GV�}�B���l:�!_YyˀtI��g���k��X�A�3޸p~��s��&}(@NB+{0A�آ�G�!�������W�$9Pʙ(EK����U�q&�F��D?T�D���ACMv�$�Ai�\6]	�Iɷ��貶�� �ѣ4t�Y��g��0?�|�L�?ͷX�ݦ`>����CW��o;������6��&qt�1��xf=����q��_�d*����}%M�'�^�IS��Y��7[�o�ia�ݜ�d��^�Y�w�SLr>s�ڇ��ʗ��U9ԉ���>f�6�[O�;�Q�;��{n��=�[���ks5�YG(�$��!U0`
}��/9X�G��Q��8�b~�p!�����n������C8?<ypև�y��w�4&oP�I�9����|�)�g��CT�P�z�}�Ĵ�qS���>�[�,Ҍ�Cog�\7�A�M�j2N	��5 �Hĝ.��H-�Ij��UWSι��xNH���� �)C�E ;f}��Y�-b�3�5�����
�����g/��I8�ᒺ\���r#_a��w���{ �[�v�_O J>A�Y�9Q���P�#�KV�j����q6OB��_�a�瀞�~���r��.{@_�W����r:���T��V�Fo[�;ޠ�^����zx��)����`�2�|jj�AbQp�O3�VSa�M���l�Ӧ·N��K)7ˊ���ę��?wy=f��/��1�{�u�C�i�CE{�u��Rgx����䭖�?k~|����H�z��d2��Q��]ɲW�+K�>n	Ԣ�#m]$J������uՂ���(%���i _~�����_׀ڼ2�I���$��� �D���9o*����ޖZ�H��ခ����]��u������@s�ܘY���TnK�Y�ȡ��Mr� 3��4�]	T-�j��p�P_'yf���R ��N��W�o�u���Ӟ�@��+sc�)Ǝ�ߋm y�l�SJSh#Q�u
!���$�_6J��:f0�^i�]��+'�"��
� �ӧ}�/=U�>�껩g�g����]ْ�!�	���ֽ	�j)��w�+��蛕 �WU��3A�4�����A@+$!̐���J�IO%q�K[�?�v����̳N˪��F̻	H��D�)&J�}�k����|D�0����Lύ1c-1鲫v���;�~�Mi\�{l/�߃]rs�,�s��r�5�!1i��eB`��{�{�٠���Vl���7���$!����XU߈Ճ���S`���XhH����j���k��<zU[�|G�}u�;��SQg-����M�o
']��<��!�nL��y=��K��艌��R�T{C��R�P+ R5k#���7~��1S������*5d��'~�6���3��G �pN�H�S��R~�x�N�zf�����S:qh}|��猵�S�8��nU|�:�P(M�/�u�ޙ���	8�v,����q��_h�x��Ťc��[���j%5��9�nn����	L)��L�Q{�+4��kc�~���,�>����2�����(4x���j���jh�?�DU;��H���o�%'La����^s�s��C͚�_�E�q�?1�N03��`|d�x�C�eC�7��#0Y�����D]��dh�B�8�^�7Û�'������U"�ʷ�(��("��'�&L�{w���D����O��n����|�C���npG�m��EW��l�����U#(Ȝ0��
��L�w?�E�1�#Y�x;FPQq�z��}A3X���=6�v�\4$�@,3��?��c�����WF��C�2�	�#�b����b\;����{�KKq:��Z�l�8�/>;'|:1�b��������}()u4[j;�^�ݟK��V,����-��6䄜faQ��3�~=�G��9��?�( �e#B9.��p�8����>��a��j��3G���Y)��+�=E6y!�E1L�Kپ�揓�\`/
b�?,\�5q�E���4����
7�*���]˪e �;���(cb����d��s#z��Y=�`O�!�`���pS k���̸^�x�����	�A�B�d�2ְ�F���~c��Em�M��{�s�!��$�bv����R>����~hs/�rY6�j�M����q��'�g k�R��K]�9��;��|$�i{��w��L���=1p�)����}w	�Ъ�HZ�2�['�l�&*��b�-+���d�i {&
�ɒ�LhPf����v��qҺ&"iGt�_8el�M�`w��Ѷe��>� T_"�^w�jcz$����=k��;���э��_�B��}A�z�}��t���˯�2�깦��]	w`��u��'	Q7{Ē�g���fJ-lB���9.iU�l2ng��ÈRb� 
KN/��0�>����w]�5�=�4�P�A��U�`6����"���T��[.�9�<�_*!#V�����Ɉo4zlѭ�C\��oD� �P����߽̈T<Xr�j~dbE�O�{_N��V�62�@�a�`�.+��bĬx�J@�"Ϫ�oOO/�̧�_!��c��!�qsi��3�l�Fp�t���{�sg`��������є��@�L���e�)�����ح*/��@4ا�[P2^r�����{���#�S�f�����A�E���Ŵ� 0*z_�k^Jm2g�N�R6v��2�ȭ7� �cg,y�����~h�Y�yB0������Ϲ��ȍ�<�⏌���·AZ����'�	L$ �k�Ғ��q��$�!p�����-P��G�sn�6�_��l�0m���lp#�9=�cW�?�7����9����U˔����3+]+g�P�i8`�,8�P��l%���@ܞ���+ǌ��so����g��F��w82}}�5T�&B���
^7��n%�:�'�Fa���YL�Au�Q\�7���(��L���/S���t��#�HX�ⴁ��̸�Fp�0������sem��	�X�}N�KE=�f�D��q�.=S_ܝC^�DO��AOB���~�[�>����F`Ê�*A�'�%�!��T�F��|&����'05c�x��������g`�a��qz�_��Rw&�����!��cB����
��*R�72m��(
�����$,���ӵ|0/�I�����k5�ì钼zE�TDW�	�\6���/�;���܆���D��+�h�X���"?'WcX����}A'Mh�D8�`��1�|��q��4�r����n7{��*`f�l�{��On��7[�	}��Juq}����{t���e�o�f�E݋�se�!w�ה2���-�8,QwiA��X��O0��-޷�b�bmw�"�!_t��3�L� P�Ϣ9Lg��.Ȳ�0�CO55T�|1�>.h"q��Z��P\��5����Gq�"%����38A��i�X�
�6�D��,6^�Y�	�!��Ï2�P�;p齵g0$2��=�VB�m�X,Ɓ�ΰ�C*H�����lϨA�U���a�&} ��?����k�8S�{�#��|��P����v<�ku9�W��y�Vs��js*Ȑ2-�deex.aBc��k����8���!�Z��ٞ�$�"�G���<��
��u����\5�P)��RH����_:$h�v���F s	�\�h�>z����K?���v��,f����4�+}o��
�o���D��d~���#�g��n��ey*�\o�����ތV΋�ӹ�L"d7l>�F���uu$(3��S��Np������Q���� K���mý���5"�����9��h����N�B��7��gk����1�[��|�3�g_��חg����C6Tq�qDY�z�X�:S�@��`��D�R=��`f��}$3C��3m�F2C���-�mUh���됱���3���a�V/�/����Q�c\׺X���{���)֤�������.r�fc)2Q5[.�|�)F�6�e��ִn��P�y��(	���������ي4�-�Ǯ��Aq�m�'=c������a�Z���mr��#���Mxb=sK��$�Ws+#�Vf���.k�"V��?�2
��.z��U8�[A���^+c��o�1�2�oᚖ�v|T�X�C����I'�� � B5��;�>.���nd�[z��z��&s�u������X��z��~�}Y!�����Y�7�PG�#�����4�4p0���g�1���>�ۤ.��E�Pd��Q��	��2�W�sS���ˡ�N���4�R���"�|�E���Ҥ��A��.�(�=�-����7��06�uS��
Q�׶	Bq'��"^�M��hC����1��I��(T�G�쌃�zf9LS�z� x+ӲEv����Ln��￹�'�a9;����+�A�ej�ӥt.���K�Q!��%��Y�����/g��c����W1	��&�T)&M�T�+�@�ש{���Նk�J�T�؋eIC�*4�Q�Ŀ�s{Ӗ���[��<��tc�[d�e�L#��j�cH�t2M9|Is����z���y��6�Y�1xH�b�y�l{}������		���k$�H��n9��6�U�?Pcs�����`�g^�8I�I���3�h5H���ԋ�G�0�*�á���P�e�ŧ�#��(�9�����1�ޙ��#���$4u��WZ>�ң���d��Z8�0ۈm��ʓ*��~���>7���tz@��wW����^����{���x2�Z"��Lbg�~�}L��l�b�&���H�FҨ_2��u��}2e�5�)Լ��� .�SX�m�Lώ�g�s(�S��\��? w���*l���4a��Q��f��	�g�l�{�xu�ZY�I��u��֠zBB��3�(��E�kLd}�С���@�D���2C��H��=jLu'�Ms�a�ț���N]�<\�e?ʕM�*�J�jrxB���X������w��DK�9*x1 \�e�m�D'荫�#v���Pu,�[��y���BY ��0��pV�Nw�Qp�Н���ҷ�+�����4^xzFgvV�|u�P֎#��J�ܸ��\��z��<ǂŷ]Lm�$Rj���_�갡�,)����F�~p���g{�����M4�5p�,џ���
#���