��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ� �t;l�������*'�հ��6[pa_�yu�����g/�U.)%��	�#e�g;�(�Y��}c�lV*�n��s4�y��a@<S���9��iwT
���`��@��_����P����iu�￣/��[��E�U��(+�X��H�\/�k �B�ǖ!��X�ܶev�J���FU{���|�W��{i�>���]�6� �� (��?/ ��C�}���-n5��r�h}�dj] cv
 '�4A��ʐ�� ��Yg$�Ƹ�˹+�KLy_�( :����0���f�?���R4��W�<M@AFala��ӆl���[�7?E	�#�0A�'͔�B!mr�j�#��wt5
TO(BT�,��`�7T<XP�oH������`�x�OM�d�\��}.hSi�#��	��<�IeD{�!WGщ�+�� �`�[��iG6���7�I��(�8y_qŤt�҂9W�&'�N��n��M��y-�TL{��	+�R|����Bͷ}���ݐ
E�]��"��^��۰�F�h{�|\�����>��@�G:����Մ!��x�#"ԧ&^i��%n�#��tȟ�5ˏ]~pW?�<ګ�'r5�՞�������FaF�"���3�#M�����:��o��X�%:DK��� �d|�>���$.�@�g�����x �D�hD�EI����eTf�X���y��.�]������J�7P�깂�G#�� WN��h�Ob��$����I�fm,1��m�rpQj�G~yn�6�C��� /ܻ���:n5\�9�ث���T�6ZX��e�͘�� awǛ��z5t��&�r�g�f�C���pJ^�?�����p��:7!�2鸑Ǝ�ǵ���`;3e�ͦ׬ʭw�j��+V���<�k�%5��.���J�2s�]6a��и^���b�cG�.}fK-�<˭ƹ:����ѕ�#	<-K5<��	�
��7�y-@Ap �|n���n��)	����%�u_��d3M�Vn�@�@��̔p�ǆ�|�b�37m����&<�;kR�_I�WF� �4����vq@4O�7�3I�D}4n�p"����?ݺ~~&H~l�(���R�
��%��hM�Ⓐ�9�4��Z4	��x����hN�f�^���c�Y?960�t�ĺ���肄�!�"K]�g|ֽ6�j�mc��&�T˄b��t�*v�1��.!�ut��ݒ''J�Z˻�[�jr��=���������H���=������@@���BD$�"���MS�6Փ��5��%���3(NZİ����u�A���꛾��a]�]ǝ��p�`J�<LU9�R�����]01�b���\�,V��VN�"�ٱQ玮�5�wM:�����Ei�&��Ir�/����}��'����5� ����zy��մ�'D��T�v���<ك���n�,E2��A=���f΂��PkT%����VR�C*Zg���:�ˍj���P{���5�eM'�>��7�f���[V���4h a��$�^&��}��������hƤehJ^|�cӠ[I�-��Ͳ]w*�=6](V�~#�!Ad�3W�(BA�����c7�2]�� p;����m�u�v��D���RN��<"z�<��F�j/a��T�'�#|�v�i�-R!���Eɞ������Q��I�U�8i��1�a;��)�8���S�e�Zh� �+#,��o��vX}�ȹ
S���X �*�X�����0\ݳ.\��^W`�+��U���y�mv��D��|N��yl����j&��=�گaX���aiP���U��=z�M.^�u��i���z��tTz���b��MR#��/9�:�5����n?)�9��A��H�3�����ijO �̚�)Y��܆�0�^�Q���}H���.�L�w���lR�8*!D-Y��6�����9��v��Y�Ƕ�g��y4S�����w������jC�a��W�F:44�YM�p�'A�k���`�}�
w��,�iOF�0���4e�U���{�Q��30�?/��Q�&e�""�}�a��E�*�g�=�F���s�k)p�r�,e*C���+��||����m�<���6P6iC-G��^bM�R!Hb�.�M��I�����^6��u��ڋSS+���Hݰw��R�J�ӌz���/i�+W'�|�ʍ��
~?�~'Ay͛/7d�	��0�A�����>�֦���M����0w{#R�=�1f���[]ԣ5'T���*#������jTn�a[�{9Q��m���jY�,��ކ8&e�{S�E+��ǚ����Ci�c�^�N�ɗU�r4Jc���7�&ٍ��
�܅�Lp"�P�ԠqZ�ؽx��q$�0����/�0>3�2���;a�¸���"p�~^�,���)TQdԜ�b�fV�m�^��L�gB��bͬ�~0g����������t�	��6~��`gI��e��ݯ�r�OjH4D+wQ�\5�%,����`uX�k�&"��H� 7��5Eub����#�&�x����F$��k�1x�r6H�݀]Q�.kz�B�tȆ��� n(LR0V{@��~��L�v�%7�H8fApg�1�����~56IШWtyDZ#"�fu�����YV؞S����|C�'��q���45�2l7��~:�Qa��g贞�2 ��������N=�VA> ���/}n��g�tW�lE-���H�� L���_n	|4x�loA6����ޛ�
;.V;�z}�̰dĘ2:��-������g���zx�F�SͳS����-	�N� ��-z3l5�	7�^�x1M�r�u��"YR�%�s�L���S�o�ۭ�.Y��d��M�{��e��A_�<�]��"�[��p��+����ڃ�͗i\�6�xP:{�p�G\{�/���!���e���~h}�]���&������_c��}*?�P�Am�t������M�HRz'�Yl�0��#5���RW���m�N.��"�����/���N�6�Ck�M!�����lbY;�֙�+�dqـ�n�F��?��c8`~ٲ+}��1���=k���U�ca�G�.���0� f��=���9�i':)!��>
�n��E�<�yJ;��^��\*�+#V�]KA8D�M�2=�Gޕ��t�n�#.uG7���axF���z�%���n�������k��m�׉��4[u=��e���!QXf�~u�Mf��N��O1���I%t������V1�>�e�:����x;��ૡ��K�f���öw2	_\��g�e�j�;K�M1ˋ6�	C�� U6����� 42M�lvx<����L9��������&�&N�W~�o�,�5��#v�[�?�˙�!�n�+�+D�ϯ���C��1�JH�<=]AW�Ԣ��%���� �Ng0z{7W@�Sϩ���K
2��B��i���=�����9�е���1����\9>AA[�q���aW�i�u\3%tY<�1�a���e���]��,���������	[�I	����YU#�%b�'�C���ͮ�t�����ŉh�6��+�Z��A�HѪ���]��#[%�i�/u�l�}�����9p6�XNr��b�1� B�hUP��o�k	S�π/j9d��|_/�!�E�4�o�{-��P�[�b ��(u�:�
N�0�#�L$���֪����`����f�H�	��{��Ss���}XP�&'����B�:�zZl�ք�,>��~��!f��,e�|JN%'x.O��rD���*pK9�� �-
���v���]'�>�-����0�_:DL�^���s�	�m�|0���
�+ͫ�kQq���M��P�v��G��D�AνgW�Օ�s9���=�����#yZUz&�w�<W�Z�~�-�h2�����K�2����7��sɝ?�::T�_����#�_�ދ����D�:2cq�o�k�}u�*V�k�����Qm*م{�!hg���9��s ?�-zd��`�L���eo�[�t�^��%�"3[�z\M��7��5P��GO��F���!"Z�J�i�v�f3E\�yL0~��i|"�s�L=!`x���$P�2�Gf�~�E;��C����đ+��R�:I�B�+�Cr��]��=�(����w$G{���d�>��Rim(�r�˞S� �@�䉯^�t|���Q���d��c�(%�ՁV�nh�6�����0�\-!�h��?�׏���N����!`�����"- ����$��l�d�0��W* �u'�G���ЄxZ��'�"B|BN;�7��f����l�;%�����ؕ�ka���<�*d�`��B׿�/���F�c2>�~�Y���͗��|`
뚊�����k����=֋�IʤR��_��)r��Q@��x��u�<��`|����cx#������E?2����)~��N���6ĔuN��d��}�yg�&�^�M2n
ϏP��q \�(�9t6A��Jܜ���In������8)�+�</��'��*�@l�
���e���Z�� -�+��x���Th#�K.m�&���G���t��gVlg�6��ʅ��D,���G�F��Q�t�9�uсpsU���֩_���b��!n�(8豲5A��4x����0�eQh��e�c�R�9�Q��������CK9Z���H�G��vD��������!���C�t��{�y[q]ά.�+�4W�y��,���*JG�k6 ���xL��_c۝����0j�;��t��_�p�l���+e��#��w�K�Z?R��Oo���a/+�n<PK |D"c~��"	�8�p�LM�&�Gc�Z����eŏx�-���d��?�V�'���0��:��A#�Խ�)#u(6��������Ӝ��V��{|�'�������]��6�8)Ǔ{���g[bN������E��lI�>����)����#��[��5����|i���n�1��"�ƪ��l��a�ɢ�P�'�z��%�	Ŷ9.tEm?f:�UYҲ��|���@��zvN �Z�>�l����	s�+�Q�T��M�lfu	�h�Y��)|��/P��ـ�WR���/�c`I9#G�|�>�y|E:/�>���֏!��d��r���X�jYvp�
��/�.�,ކ_$��5hu/\~��x
�
y9+2�/��%ɭ�5;�4=�s�pF�n�_�d4^yW�F�Q����k�>�Lػ�p���
��27F�MJuAp0�wh]fm-ϓ NFHWfY��1�jD������\���iK��9<T�ѹU��-y�R��뷌aA��X&R7Jf�
5;�݌�zmM�]w??�MT�=P�{N�}�"�B�C/�X{�ҤH����v2kD�U��������KJ9��K^Hָ�m�h�؋���c��*}+Z�-�;6��B5#�S5�u5���6	(ڒE���Y¤fs�舡0�EiK���#�q�Ћ�� ��^Y5�c� S�!>D�m-ɉ��&�j�$S| Lu�m�ۓ�Ȁ� 糵>��$�2���Ku`���
�����0mR~3�p�eQT|���u�wz����H8�m�9�*�r�f���GƑ��,�u�v�!�o�1b�ᱭ��Pd��=*����b. ��GI/ō#s6�
��X��#��.S��)��q�A�@p�L7�8e<�R"��Fx�l�Va�W$úM�݀�t�Wk"M����u�ƀ�Ra�L3��\QS��2&�tZ�V�� $�`@��OZ�;<��;័f2�T��W�&��5�r�m��	~�ޝv�w�ts��/�$�k�[y��T��%����G�����="��fӰ�Նc(y�����RF�)g�����c���i�u��1��d���TɘK�)9h�x8����[���n��Rkw3a�i��q�K'I��Q~h;D!���!!��P��zI�CWmD�
vYhIXꜥ�D>UA���������_50��9_�y�H58b���R���+��0�X������:��QlI�O��c��4���7��.g�_˒����G��h��H	<�镈�7*�d��K)��v�7{�dcn5�;R0�	u�m�/��E��D;�9[{´�ߨ5D�`�RM�7�]c{%�j֜�w�߼�.��	<��&H|����}�Gp��D��T��\\�D<����Z�@���C.��� 5E��tp�\3�O���
�hB�6Kџ���m"�a�]�zZ���hA�I���1��/V=�ڠs��Ɋe{`\�NA���i�~�k"Bm��٥c��!�ɥX)�ԛ~4%�����U��Tu�?����r�}iK��D�t��3'����N��	:e��A_'s���u�c�)���-�'�*�tx�bꄘ�ݯ1p���[7kap������6z�%�0����2Ȭ�.��6ƇH
TC#�s��<���}5��tn���0� ���2l�<�uAiعK?�^����㱷b�7�� Z}��T�3�-S�[�v��/=t�_�
ry=У�o�!���З�{�~����XD.B��/���-Y�������Z�r��R(�y��1ڡ����C�梽��*���V_?�:
��<1�'8Z�������i���FY�ԛYЪ{0��Kl.ː�ז��g��xߤALE{�ɲ���	4�з~|�
?���,y�X�tX]N��l��i˟'���5-=����$�Q�TZ���;��3�����u"H�P�0��T��o�Sy�W<����z:�/(�ہ���>����N)��R0��?ndu>/#k�G����ɚ�
��s�D�%w��E����/���*+��K}�d3�j�>
�m}��!�Me�A�qH�@j��h��@�B�R��m�+�@"�H���㦇��<d�9�fLs�Ep��U�����.7����&�kx�a��y�V
$����
��������{3�s�/���I{�8�hyіk�����q�L�+���C��_��֎7��+|y�P�	ks��20����Z��1h��%�i�͸�׭M�W��"h�!���>�Nrs`�J��������$V@v��� V�Ɔ<E4�iiZ�M]�����sG����B��2���۠���G��s��M�=�m�z�'�(V�<_+�,���G�.up`R�Jɮ=��$�z렜�$7���[�	��e�ث�͢�ǥ��~���۪gӦZ{�,P��ΪPb����~e�2V�
v	�1�-�b�*�,�F=mS�|#�]�$��LB�*�*�?�T��JgfV�%�%,�X>�����u�
<�j&F���M`��g�ؐ��%���9:~`S��5E�'���&�ۉv�(��;��1O�x�ګ���a�`܏�}z�����SleH��o��,a�!���b}�	�_�zV�dO][Q{�aa0TF��t=G�E����E4l���A�`�񺢐����i�}W�{m�s����k�a3"��e�wE8�9+��,����nǩa����t�D�����)��� ��i��}
�(���Q�RUK�e�)���I*vB�O��	Ю�ģ�tuؒ���\ I�<�IT�,,X½�F�3,�
�"�sKs�ļ�+�2EP�̋����=�)R.�<����)l*Q�C�������{�r�0�0J��s:b�~}X;~���#�I����EPh���+�.3�=x	�k1,�b�.{`�UL;�Z�a�g>������A�!6��Dv]+?�s����D]~^۝�V9�1-S7���`������r㖫ژ&{�>�{�d�V�f��-pw.��� N8���d����Ś�<���7�i��,ax�� �iL�,�5�Y�	�k魬���ZVU������؍�ͷV��7lF���Gҗ��>�"B��h֦���+���g�:�׻�\�B���v#h��V�
� �#O�2b:#s�r p��Ym��k�(��?ZT��܁	���}��S�<�qV�*��=+Q?����S���_X$���)��J���?(���k�L��g�ɯ���Յ�?=&�<o�#�DB(R9��3?��}�Bf�{���!�3�VR�H��g�&��Y�nT���b�!���7���|`X�oz���C.���3F��{�/ӛ�"ے8�E��ٴ#���\_��.���;�\w:;���c�������n=�*܀��S�����Zv�,�y�I���:��su��}�N�bk���_M�^#�x;�{ĳ%z�3#�����%Y�מvE��Cs��d0Y�� "Ʀ@��y��>��k��Q�(k�T�eVϿ\S6�tK��]a���� $oz+�t�6�򑋼v��f��� ���W=�4658n�M�pn>�-'3ڦ��H��a)}l�<�k�ﾖ	/�.K|J�0��@�5dbT�:��a�IE�vO�7zc������C#�h�A��r$�K��}�⾧���	EW0ǿm�t��!H�7uu���
�'VP��$�u�(�E�n�a/�y��^�<��hȾ_;��8��=����I�[\J��23�7�9�e�Z�z��o2Fk(��}�)(�Ϗ�k�b�g䲒4�e��K���yo#��mM�^6��{$5}�Mi-�i������)�c�|ޤ9��n+�a^��6�+�HUp�W�T&�n���_�G����'�}cL��ғ@K8A�'�cw��(����"�������mfB�7�[~�E�^��"V�˿kL��W�T��I��&t�brP�˄5��Ѡ@\���J����s:�f�N>!���ma�#a<�n-�F��:�z�[��T�o�=0�@Q7K��o�܎�	�=5�.�,�U)�WU:����|6qP���~��4R1V����[�0�5���t����La%�샖�P�[�}�i��v�ZI��mZ�݁���'�؆ayk�CV����~���4f�	�4̧�A�4�vSlH�޴b���/���x��-q�
��mA�ElܛB9�Y�_+��_�jT�g�Q�ؤVY�"�b�,�s&7�4���[U�:�����h��<Oe�]��a �₤m��p�����������-���X��.�lt>�c��x����no;^�n�?��Ͼ@k0�����:�9� �C�GA��/�ՀU9�t�TȵI�9��'����~&>q���g� �"�MF}�{Y���U�H�K�.�q(6�]K���8��lv
T�BB���@�=O`9��q�]���&1��f����,|�C�!R���ґ�;�9�ȑ����2���N��<C�*�j��ђ�{rQ�CP�z���y�W^��]��0��N�a;;��i����ٺӍ%h�9R�cy�!�Yh�O��p���r�z�$�C�W퓚j���2hU����v�v�%���Y�$���G7��į�i�3p�Ej&ߔ �j�'A`r���$�n�PJ�x�{B.vE;"��>x�CYu������7�n�l�~�J2l�6�L7[�_��Yv��X�5yoL���.��/o .Ap��[���i�O���ד����cTZ~D/qK2I�9�9���\��d��f,�r�-F���Ȩ�ٽ���K~�s�L���8[�����vv�!-Z��?ua�2��Ȣ� gg�=~D$v���F2#o��*a(��Mm��y�h��|�������%Ag�x�����}�a�XY���3gM`���QK�(���� �(�B�f8%�ٶ)�;:��EN�uC��i�%��-����#�7�i�CE1C�$`5F�aI:�.=B�nX�U�V���D�+������?�t�LR<� 4�r��af'Y
̲L�39���rOP�B��Ҩ�1v����j�9��m��*2���N�Gs���nh��r���Ym�Jz��L��� p�S�_�P�<[�t�f��A�k oT!�����awn#60�[~�2o��"_�bh�04�����nα�r��M��5��T7���)$�mIK�聤b
�ْC@Y*�be��c�dijJ��ǏZ�����t�);<,o�B���-�wLs�	3�@� �(�fI�{6�1P�;2�n���"rF]�� ��LؼׁiS����@8٩����N�{������L�y��+6^�ʔ�=%Wm&Q�;"ޔQjt���{ILH�l�ҕ���W��p�=]�w�a>���8QLq.ּ�&��,=��a�S��t��+����=b���<�2C�q��`$�'�)䫌=m.���-I��H|Z+$'���pLX��
�@�鰼~*��%~������L}3�����-�����;Q�D�&},a-|�����VR,�WZ�(~�[��f�����0���BT�۟�"ѩvo�?�!U��D�xw=@�{o��
���"R�����5,B�%F�-��cJ�F�3"�r��D ��=T��5�flG��jJC!/E���O�*)j��̖N �Z&���|�,PZ��u�>���x$Y�����<�� %���^��K:G��^̌�ZOؗ��9�U�+Ie�s�<�*�d	��T��tj�?Q��;��X�N%,H�KNK�b��Zqҙ6����t�~���b�x�Ͳ��^W�R5�%U�rǗY��j�q�f��b[䌣�����/+�f�7զŮ�1��������T+R�v�i���n��EM�衚ڒ4:(�p��5TZ e]�2fK��T�@�*���+B@\�v���2^���Ƹ@^��Mc�5�C1�8S�����7T��@�UX4џˡGL��(����i��ޖ>.�r!!C��d��(#
O�p�X���l��˔������D��,���
)Wc�� <Ry��������_
&Ts�w����@a]��u��m�P�x������g}A�:�癜Õi*�篸p(J��ů֢���п�>��+��'<�U���!��_Y
�ԇ�tr+q�F�@Z�_Q�4�i��F� ������"�h� �h< QQ���tW��?�?�X9y�n���w{\��P,�|�3&�TY,��$�������"��n����I��� ![Rw�:_I�[�pn�����9�3rD�@^�4�P�k�>���+{�0e�J��V�'L�� h�8y1����ݠ�xx|HϰԜ���=�,�y
3�UЋ,�Ե#o�Բ�_p`�����
��NWz!ا��̧�p�-���/�n˒ޭ'P�1.��j.���ږž�.��M�,q<��e味�	k.��0���[�JO$���*}i]��Z��N� 6d����1� � o6K�+�ګx�R<��>����فW�ضA֫����WA2��j�k}��Vz1+���dmn:L�K��UG�\a���gjw�v�P]-�6!!��i}�~�*}-�H���j���tIP\���:�/g�x��@Y�Ȝv���ĵK��`��<����F)({�N@��}����6�`�����5F���!�5#Q&R�	�q�)p���vH��_�bݿ"����L/ Wpf��0�ŕy��nO�
Ϊ����L�^֮˘�}� �^&vA1L?������g� f��bN����|N2G휏���htI�V�G�=e���WV���p:���_&�f#��,��&���' ud����w�_���:䱹ļ�OJ
��uS�6��G2c�����o{�@�LU�(�|�s�߬���s��Z�+cL���by���&�4����-���{P�3��M�~mf#0��=׌|��X�O��m�f)�´��gZ��6�L�t"@�s?$8�e1!U8a};�r%AA�c�w}��N����o|��K
~~Q�Gt�_*��ȀTN�:��#�?�݃�l��}�k�Mtչ�-����L���f���i9�����̰U���S����'���M��-K�F�a{��T�H��V*�U��i;������_p)N�����X|�5�S�4��VsC��$P�P��Z�!�qH���?�I����"X��/�΁��s]n�K��;�N�fa�B.?�4�0�B;�4"�2�L����tr���X!�ņ�We9\���,pg��K�gi�M�p���Qٗg2)z�;��ѓɞoN��lk�Xǰ�_��^H�ह�w��	�1#���c�W�(��EM�Ň��$��(�:�,\��A}IU�X����~���}�� �Ҩ�E`Ϙ����,�|�mƒ��� jݤ���-���JEy4�t%�<��;,Z>
	��2
�@�4�P�F|ێ�I�#�{>�~��'�c��v���͗1"����P�w��͞���{-/�\`׼�j&j&�K���$Xձ�k�l�+k�Mm�C�m;) �r��?���18`�Z%$�q>��0�EI��NSTS8�X����b�����RYe"���Ap�Ivgֶۢ>�}*��Ѱ'���r�f-�ÝMUV髏��~&��=@p1c6��B���X��1��Lu�T8�C+C�-j������J�w��X��_�)d�~�ՂW<�� �"fo�t�`�9@/�"D�K�W 3�Z!�~�ƈ��w���I4e��$0uK�<t��v����-���Δ�	Wn�	��3�}��N��~Fi����`F��\3@��
��<�&c:��HW����E(�l�8����S	${W���e�������z�]�n��TB���U���x��޾����Hgp�7�;Jza�On6��<T�]_������z�nea���;�z�%�R�������ee�:]�j�)4�nq���G�2X�ѐ����ċ��_�������V��8�R�'\�����_\Jy}��ڋ:ܗ1cmEf�7JꆤA;aV�;�_%��_ڻ����TY:���6ā�tg������J��3G`����@V�%U�9�kkF�����tё�5-��G��H��l���?&d,%JޭF�le"[����y��̍Nqb&�2��9�B�.��m�3t��=�uA˥Amp#�{ǅʱ�]r�s��%�2����謃+�>�,�Ճ��2��>���s�\�[��+[�ᇑj������n����V�P}=���7��R#!�7�}*v�3��ӹE	�_<k�o��������ݎo���0�p���?�}�H8�c��$FYa9(�8S���V����x���B�ܵr���{t/��Z�\�����pۆX=��~��Ʒ�7fQ7��[>�,���"P,�7W��<O��iL$��+��̽D����\�a>��4W1J0<ImD+�
������&��<84�N�̣��˲��[�%��!�w;\��Z9����n$p���G�5��#�]���P������s�����=U^�Ի��\w�g����.S�	�m�#e�!D�=�Aޡ��U��A ����o�H$b@CL�=�?���]��j��bE��:"��E|��u�e9��]�XM>X�d*�~:gKI���媷}li�h��Щ��܏*�.Ma�V���)"�X�L�J_��,ʶ�C&�����	�C�|u�+�o ���h��q ւ!z�mi��#����o�k��-:&ir�&w�C�����0��N9��V����e�m�=l�a�*Z-���Cl�� z�2Q�NRm��l�"W�m��O����Ƞ�5����T��PAY�d�1��x�R�>R���e�md_�~N��֯uJ�;�_4Wo������_H�A�:��Y�W5�r�B�jрv������D(�\-F5I���![���#����5������ɽn�Ej�O60�~��Rߨ�H�4��^t��¿�Ƈs��j� w�6���hH@s����2E�܎q��ֆ�g���;6�$�Y Rs��`[_�턾�w����~�~����x����J�U���g�rt�8�7�'+��P�j���[���ҝx1�7�{�h@����O�[7%� a�@TRg�;�Y���� ,4�g�^���:Z��H�nC���Sެ�%=(+�A�9������t�j�󰾖��ʐ�Ǝ�l�"�N��t����Z�%')��¬���l�d��鋓��t�g������Z��䎰�s�y�M�.;�J��j,���?��z���ߊՐ�� �4m ��p\�KA�r�*�V(�'��O���Ĝu4u�u_>FsV��Q���ortWݼq/�xO�)�����(�k���HJ�U��.�	)@X?º��l������´��Z����,�~��m��M"ɀc���;1�Ѐ#fюb��AE�x�m�%�Ʒ&�2OI�R��)���$��=�N��W#s��,<��Q�a��B�`�����'P�`" IRx�p'R\~B���ٚ�p�����-�eS�&W���k��Dwc�a�Z��j��;��SAM�Ԑ�cpN���,��n"�b�_F���M-0��Da�q���#���L���.��A�cl���G�bO�z�aᚪ����z;6�o�d|M�=�z�G�q�����v���j�-��D�(�@����\�.�S����`��=�7�LS��s~���ﰪY����K����\���a޿�VdK��t���I��w�N�ݟה�X�_�=�8�|����<��Y �3� �����Z��桉�) ax��6�;l�%z�1�����O���5�qgF�y�cѭ�e[n�ɤ]n���(02�xg��f�	>��F��h|.��tf	�3DT\�`�Z��i�����5>�3������>�Ǌ�_�7�d^���=CL��N�?�c�3gf�9�OD\���-RUy������~)��H�<��
���h"�Ĳ�\���X��mO�[�[���o�/�%&	rL�$��C8I������]�6&5�\1p�VtX?�°��ۧf����b�}i q�����<N���~)��I�in�nu�P
��
5��،����;G�R�\]H��7�p~94nk����74UkF���	��_�$ �$'5��#�f���n!�>�ا'�u4u�ҵa~�����G���hd���l&e��W݃���]��{�X��Roz`�\��0?��Óg6җ-����`�ji��
�Z��x� �4B�&]�a/�J�u!?l����|}I��y���U�p��n@P@�5j�F�o���^���(�l 4Cv����^�z�^v��YT9�?�J��黔7G�- ��j��!�niU�a?�J�j�0P[Ј>�ߞX��x0�R:E~`���v�,1x���4��KӐ\i��f�u�Y�P`��\1�L,-B<*�;]��ٜ���mKqڄ�3F����\�>[xF�9Z�|$���-�����F�qvT�ڏC��l�h�E$�;w;Ŋ�%~F8)�;!s/�0�
q���|\��}��Id�׋?��8��K8	���Fo��Փ`�����b���Є��=ҩyI#%|o/W1��J@�d�ԁ�vk�b���0"��|��S����A�K�٫3.���@.�"��V�v�CG��1B�u�������c>0/aW�;��H*_%һ<[�������6�=C]���h�S\����>c���q�]|;��h�4*0 �[Y��ILकn�p:��S\x��L��,���%��F�p��ć��q�%X"�-��҃<bpBL���GΓ�~���\`oS���K�]x�L�7�x�����?�:�fQ�)�c^�D�\XK�;|ѱJgȱ�%���$E�-GS�ǫe=�@��Ƌcۅ6�G��b��<�~�&�][2X�8��>5�i9��7y�����0UNJǋ�ԃ�c�B�B���x�V� ��*h�F�p��q���وY@�o�JQ:�@��r�l#I%4=]�e�T�H��U���uq��Ş��LX�f�n	��g��-�MK�"椔Cɡ�XC��Û�˒I��\Q(6�l��$l6���U��a�� H�bn��d�t�{t��� e�F�\D+υ{�lE[�ѵM�th Qצ")�h���9���|���AV�3��5��'\P,s&��C�]�V�i��D�o{��ۤ����ʍԃ�/!�����4��"'<����k:��d�k�+�K��~�;42Bc<��*+�ww��ߪ�%-G�{f� (��S��d�x�#y�� ^���|�����ÞX��SS	����<-O�Yb��� ]eZ�����V~�qMG8_��R%ǿ<xv\s�w,��N��_���>k�٭���t�C��`Sq��):�����p�&±�rE+z���W�<�"��iQǼ�WPmb�"Ї��N���/�`0#	: �}���uuDh��6�JE��ű�b|=ڮޮ�����5�#�z&``��U��R��\��i_�L�g0?��h�
.�'��}IU1�X�m�`%�2�S���"��vj5�q^M�v�s��E~�$��|j� E�����\Ѹ�<�oB��WG�����u��2�����f��o��H8W����}�y}=|��"������h�V-~�Z�l^�9X��_�-s������%qdȖ�<��'�6�g�"��t�P�z�լHz#��7�_����#:����#��'q��;��_�hW]��pwGZ9&����W�"��"M\��d�4���������4,6Wo�1�xJ��?�{��*�ZT,(T
<��҄�x;���v�����9�����qՌ��E��	\U(�=�xG5	�W���pO���0Pë%7�d\��!�2�R��#�%J�RPK&{�pj�̝����4{a��g�|�߁�P*�Go���o~�A����!W�nz�oP��y�d�D��Z�7�8�/E���/���H�TPN��>��? �(=��~�0�&G��R��V�0�#�i���g\��xiο"��&�-P�ݧ�<�?0�x+3Н\����ǝ�!fZg+���̖�>[�c�U�t�p�3�"	wi(�����[�D:�����ce���k��)������')����z�uQ�ݿ��b�&n�!�&���Vl��"�c�W�o�Ga�+J�k�¶�CvC��<��|N�ݎ6l_}�M�F-�*�29̿q�;�鍔6pL��h��#7�;:�
z����0�r����D�+��Y��f�>n�"O�s�ͺ�o�E�(��oI|ڠ����,��lF�C8}զ<����M�^/F���D�B���I�n�����_�m�ݝ*-ۓ)g�_ �voJ7~&��{�EB�j�l�t8EJ>���1 =�0�\�^ޯCt�
�,��<3}C�)�L����]DHLOL�}����⧏���6�>#w@������-wQ�����=��,����^R#=hST.���n�x�|���w%4�;5��g�5\d�+��X�=��J	���ڃ���P��T:�Y���j��d�r�"mgj�1�럴��=h[}�8]�K6%�K�#|҈�(�+�@wV�C��J�8�,�T+��9��̒�倵,Yd�s4�@�G�*�q������E�m�7�W�ʑ�'�Yo������1���K�F�	�.I��I(b@��jo�ݐ���'��HO���pY�7��W����+��M��B)Cf���Y�!b���o�f����g{�U�3�:�����TJ��Th��r�(n�P5�i���U5_ē;�����UV|�UP���W�����:������6+��}`��3����G>���]��{��7O������q�b�k��Q�WiA#ܯ�����/t�U�շ�{���)Z�D$���E:=��,��^��ܠ0V_�J���VK
2�a�Q�G4�����PĔKyRVx�}B�I
$��C��s��g �U�5<�Sb��%o\�j���笖�2T�,k�=�x��`��tr|�ਂ^�d{BM�r]���+5!GI�2�^)8�ku��<���1Z�Rj����%�GuU���c�����N� F~z���BY�a����`'�iEQ�F2�F;. &����J��Oܚ6�S���*H�\d�Y�BA0�Q���Ķsr ��s���������8a8Mt|�eC����o���,&3'g��j�|�x�{$WM��j���`E��q�OFC7�(��v�&r�j�V餴�Zb�"��"�����&t������~.�^PP0W��\�/oS�-�G*��<M��X/Je����Ub���ZWT��L-���h`�$0M1P�ʠ")�ih&G�0��UmXA�+�e��0*m����d�'q��M��%/v��Q}�`��7�����6��?KK"�����}6���l�ywrp�E�%���#U��_�q�{���Y ���pu�C�0_V�l�U��[��Yi�@+����j��A��$D.�cζ������ѐ#x^�tZ����L����/{.p4�=�#J8��Q�����%S���)�;Lq�b*ʗ|H���fIR��MI�f��x��]h��l�T�_��i����?�d	��]nS���L7���� 3�RL���Ǵ� h��6����2d�R,�rr�+WR���{b�g*ٚ@-����D&_�w� ��0����(��T¢x�>Z�#�cY��z^u�
��I�D���������_)��q%1�O���̻o_.�[�gfܒ�/�1�|צ_�L9{�IOK��jp#7���P~7<��?xZ�Z0K�!�iJ�^���Y�t����m휺"3�WX:f�z~I����~Z{��I�p������ۄ���N:F5&��|���!'���J�W�	��STT��>]T��A�K�7�ۍ7��)��j�N����T�RaU� rQV���KUW'����D��C�578f��J�{'�r�1#�iJm�����HZ.�h|���2q,�X.��I�bvO.S����Rq9��dm֔�0�Kڼ-�Qr��>'�Â
��־��.�����P���\����A����!�z�'x���0���߰����Pз��%�v�I5t���v��g��L+��̅)n:�wsʈ���C��r9 β�R�n����-;q�l�Ĕk⏾���T�d�h��p~�����6��{,y����=	��D3呛�Ӈ.�(
����-I:��Ǒ�Ow>*n�ɚo*��5G�x�, ��1:Fa�Ju `��væLN�olfߡ��@��I���J5O�+1����͌�xR��+������_�n������w��=>�or�?�c��5�ZvUX�Bj���T��ѣ�{a�v$} ��Y�z �M���
i��P�����/$ls"����;#&�7�c���dυ��]�������q�[A�3Yt8ٷr�u#����+�z��������������ˤ���4 K�>�z�f��l�Q�����Xʥ�ӧ0GVj5i�X�ߡ;�����l�|};͏�s"�辔_�ok���c}HM��Xy��`�K�M1�-����U(29Q?�O��±:��r`�-��C�S�{��/���=�E<"1�X�|]�)�\jc&��-��;���\�u^ul��A��W���(�s@ʑ!��s�un�~q&M��d9B��R@ �{�_}��k(��,qa�
����᰷\��i�%�n�����h�j�{\OsL����9��<�bf0W\k��Qf��:�2'�8���߹�hA�&J��\���ըT�j7<��rOi�y�$�]P%Q+J����:a��bE��ɓ��[Z`x;5��h���Uo��du����_�)��p0�4����i<@����ߘ:�t���w���F�g�M���~n3�	|��-Kk��~A�L�l� a��s�J�`)�U;�)�s]�$�`�o�-0���Z��ڹ�[x;�~��BS��+��Ǿ���v?��	��OU/�R�c�Q��m��";2�Alo7��=�x�6��CB��@P&���h7˿n��&�>��8|��~�0z��
zد\zS�E���:}�if�����T�١��}VV�(H���8�S��?�g���2pQ��'��&~+�_T��n��!*�Bq��Bz��i߳�k��Fy9J�QE�$F�S]��:;�(�'Ycr�,��O�� jqָ��Eq����|y�rIj`�5��^�E����L�`�W�C&���Y�(k	�Ֆ_l�1���8J]���������f�nT�J~x���6 ����˥Y?��3"������.�Z���r��m��ҹC��YW2�7��_f���650m�~aݒ}��q[z^{��$�`^� �v��]H�T�n&�NU���x�^[��Fn�{�މ��Б�Ր�k Qxjp�]�Of�4-�eDt4���Q�vnfH��#��a�J�a7Xv��w#�p��G!r�@7Σ�~UɢWz0j�$�ؑ�N�=|�t�ױ��d	TsWuz�<9�H�>G��,�Z�j�Ğ���5��i�;
����wvyTs�w��X� yk�:�'T�x�5��X���������oa�k�<��8)�=���K��`�t���u�*\f�@����D�����6з�Ĺ�nP���DgJP��;;D���Q��>�F�^i
�X�-�x�S��a]���a�T�1��l��Z�HqQ̶K'r9d���mn����e�_���YRe �%A;5Ι�s�{���d]7���<AUƼ�Hq�K����W<HR���X�o��z+�DU��z���X�#�3�X{�dy��H~#�膤�=���nG�bS��L �aOq�Ѕ$:|4A��V�ey%�]��(v�4�k�ܮ��Vq�RSv��2�[v��op�Il�pRޘN����*�C��
�;l��׸C4�~�����CL��?m�nƊ��\�^��U�ZrJ���ԛ�K���,[T���*�f%>�����hV� 5��T:hV�-���	m̚��G��;.N����n�B��<��W��o�k<@�Ȓ%��w�(a�G�,�L�u�Q�����;����W��	d-�4e	��fuz׏�"��z�:�YAר|�DO�"���(�@@��@z
I�l�i��叹Vt���]ID:)��`��q�2�BU�$k��ΘFo}�mA]��R�K)�!x&�Jg���q�f�q����}S呥3|j\#|P��Tv�/�ު'�ˋ�!ubQ�Rf	�L�l�  �����ji�1�)J���Q�����	S�$~�1�|݅�h���*�r�~eG�o��T�Ǥ�aczF����Z0�&����I�CSVo�#a�d�3i�������5[x{
��|�0ZLj5\��Q��ȂA��Ǐ��i�����M�S�?l��Ԅ�?!�=Yj�g;����z���B�T�_�����}��%��"�I-����`��/��W����i 8��$xdW��{��S�����:��8J���q��j~�k5_��[�9�ρp�<."�'΂��<����#�Y�CI�|h\*�?�9�l�
>���__S�1���̾���]sBA"�;�b(7]N���4W���`,�ݿ�ܓ�?BA��Ɉ�o��"Np�1%��22x�Bh�/����W/]@H|/Uo�@�!�{έ�'͜�D���[�V���Ͷs�I��e�}��q8�&|6C�n D�y��`��ǋ�ε�@Nm�m����s����5��\vy��@�i�\g�#�a��z������b�8�|���ߗM��_HW��|����<���g����Eȯ��c6��k���x��c��^����y��Vc���8�̻`(ʨ5�S�v o<�f(�G���
�xI� 5dں�z##-�XM�Ol�\���\�ǲ�SF�6Kd�F��]'Uk��h���6X����y��J�S�R(��~����.�|��9�w���Լ��܀�y�O��J<`���7W�ö�p"�k#��������1o?7�4<�E���R�/n��؋�iAT��$���Y���.Xm�κ��Y����h���\�j��i�'J?��D���{�LȲzt��iQ�Â"J�\�Y�v��IW���=�����<r�ŋȰ ��ȟp(�Qt��
q��\{�M8�W�@>�h�\O~eS�P��'Z����6��i����\Qѡ��@F5
�K^�
ts[urjJ���Nc8E��6�YW�]"���)� Br5���2ʇ���e�4��7�
S����o����)ȼU�0�X�<���7�i��kGuҳBI���$vߙ���T��cY6)���)��D�����OgP�Pv��`H)厸T ^��|�����A��I?j4�����E �N	1繩���<��W@�R� w�rD�������X��q���gЙD&�5��|Ռy��8I]�1�V�M��r�S1���s�h����Fr;9\IL6����-w4L�|��E��ˣ��M�p�X�4()k�;`%�`���v$P�����׌L�c[^��G<J{�~`]��#Za�q���:V��X062`"lI�G0�'�� =C׵��d��ɧ!��ڔ�1(C���������Q�l/:�M�Q;{[��dﶤ&�X��~"�����XHJ�Yȡ\�<���f6+������Җ��w�^�coW����_�����'��L�=���M� ��Zګ߰��/-ތZT�"���6�[-�*�[�L� ��t�(����0���U��ʦoy:�2�_�h��:$~~/qD
���5����ɞ���+���i� F�Q�}�07�qM[�&Xjɋ��}�N�p�3�?����
��\�HD��X�xHG�lM\b�g�+^��Ar�O#g��sHae��"PS��MRɬ[��ofSFYi�mn�0PT<�Um��(�&���T�<|���!�.��� ��~G{
ߏR)�z�W��J>k~"e��8��7�V����/1԰[�����������)���vuK�Ĺ�i����������Ty��b�Q9�=���:�'	�̐)�}�H����m��M�BN:�|�P2`Q���Z8o6 ���~�@j�C��SҺ̜�(����y�i7'���=����������G��Ȳ��{�j���
8���G$��[��/O��G�c���p^�u���?��<�yeY�z�����_�c���@.e����;N�����,c6�fO^"�Mj��<I��l����n�_�`��2���t����+�|�T�6C[<��j�;p%����'�v�u�_�3n]P��Dٴ������D�t�V��qȩE�1�,���)H=�0Z�d��8��UB�E2a$���T�̾�h�q�Oa4�u=��ˑ -|�{��&ӶtKz���R�&����7�5.er���'�t�ꠤ�󓈻9M���� @��Di^b{Au�=־ZE��K��=R�x
K����	<��d��;Zvt؎1�=e&�f��e���q#�)RH�}GҖl�H \���N�K���a��a�H�#�@#�$s�@���X��ʢ�`��"�.Ş���`�+'����b��d��,�%� ap_�+�:K��U�I�c�a���7Q��B`�}QA�^1l�Nbf�Q<�g��Ўs�.��Í�����y+1!���BI���vI�!Z|tu�w�(S��)�r�$jq-���"��o�qR�*%�X[�,F���
��~xH�e_B��_C�� =@��
���k��Eߴ��غ�ĚN�U�sbk=�\����I� h�m���0�j������g����Uy��:����EN�X�P-wG����b�G&x�U���;�0�R �A�hu��O֯	W�:kkb� ���ԛ3z�ɒ������8Я�e�Z5��,����SQ��V	���7K=��$m@�aP���H�r��(�[��1�蝭����劗���OH%v+8����,�h�b��-� An����Z�v�j��M>��vdq'�i4=l0�肰�� BPD�g	R�B���Z�e�C�	!��SS�Hˮ����8�I[QX=[��K"�oE$\އ��W7z��������|-��D�.P�Ed����#1�(DH�^�_�Ĥ�^�Zq��D�7��ipKv[����Ba+����H文��h��:g�=��j���M�m��}5>�H�fh��Q^�p��Ĉ16R��y ;CYs�Y�a=`o�o[��3!����	!v����g��sfA8ӂ'���D�}��4A}!�d�c�an�Z�ie��=_`�_�x&i3�C���G,�EI��O���W�O��([��`Q�Y�Eߜ��rpm0�+���W?}B\[*��_as{�J��vC�4��q'@��� v���q�wP��v�pL��:�"���\�F���e����ˢ���_��O�w9<���z������&$��{/%�Eq�d����h����R�ѥ��要$� $1�X1��C(�3�"��!^��3���ba��]���C��E��Rl��2z�#����G�ۯ���y��WH�!>,,a���{��@����9��)��'��9�k�	>����T�����O�y%UK��Ir��`�>��Y����]�v�/�ŭC_יS��w�?�L� U>��J1z����bop��_:'�d�	�<w�n���}����櫡K��;��[=����xiK�$�ĵ�t;��,UY�=*�3��.��_����7
,����2����|-�I�[g����C���t�W��nވ^.x8]��bFhrض�f�{�N�d�)�Ҥ�� �ف�1�W��"Y|8��r�I�_�Q�,��S�];����2e���.�e��E�Ŭ�ڻ�\#<\}r@U�A���St����C;�ۻ����S</�O,NcD���E�������y��h�)�/�������,���^2B��M�M�[�ꨰ���)ă��k߮B�"���;7�eZͺ��(Sw*�C��0Rv����V�v�w�j�Bi*���Z��p+�X�]�c�<:�7v�_ѮCi� Rd��������l��1�륧�}@1�t^�3ܵ |�B��܁�ү�u���?e�R����{˂,;�q�Qb�������LX6C���ⓡ3�D���.��5�t�7����үU�~٢r�� *k��r���k��� �tT�ՂSC�NAZk���.Z�����:M�E�Ī��$Y�B��r]s����v<����E�yS���d~�g�N	�IT�ȱ[�d�(@e�{.s�ֲc~�B��$p}#"��T
d�/7��p����S�Az�z�/���6/n�ܶhu���5aJp0eE��H8���B)j8�����m�6ƞ'��=N�jSmd�2��Q��]&��L�}{ZS��E�����'X?�s���p��5څ�s�|�p���4�+���9鵿���	��$w�/�����H蘜%7��uncoЀ2��~@���T{^c��)����i�Z�p��3����q8�'q����s'GhQj���?,&B!�/�$Y4�	4"k��Hs�
���:�0��,H�}tr����#��P�W�r�x����	l�cg�i��a9�,���J'�ikƦ�֨�3F���>T��zD���7Q0?	5�ji�'_�.��e�FD����:�t�|��/V2z{��湎�3�{j�g� 8m�a$����9*��*凜���Λag��F���R�Nq/ں��ɒ�Q��p�Fv[��z�z�z�*.z�_���_J5�\��Ul���-r�z]��#҉�J9�P����&o����x�sq&p.�-��pF����}+X#�;���gA�Η��Y\ͣ�Gy�`��7�sz	��m)�-]�g����� W�ot�F�/\ü��P�\�V�*���z\������b���L^ǲq5����|�F��Ny%��?��#�lE�n�x�> ��5`�J\U'�\�*�<�YP֘y�.�C3�x�00��T�]��
aTvM T����SY1�Xj��
m���Fv&A�X�������Fh[�0��M[k�ҍ>���b�*��a���S������&DtC�X�çυ�\�@MOuo(����l��Љ�.�Jº,�s:���49살������D����K�2;��3d(��s�H��ޘ�A��m�������m��52/�Nڒ��g�S��B0L��3��f��<�ެ� u���>��5#\�>z���:�gg<�'}}�썔�L�^�?�π���7qJ��?F��)lz�m�?�Il2�ZL�{����tPC.i腡�xd&ϯ.�?����GQF�T(�#�E���ܹ���c֏'!fO
�,���6��S��퀔�=m��E�p�?2D�C>�`��2�D�IQ)J����]NI��2h��O4fK�V�wΓ
;��!>:�ũ'��qp���җ�2�[Xw6+�8KǬ��"��C�E�"\��TjD�mx^�#�����Y�߈ۂ3Z�g�l��5Z�G	�:	c�ρT����p%&-V���ej �������h2��9�� !�����ˀ�����X�3���j���PA��p�ezصd��j��۫Y��H;`�E��� ���A���7�W߆�S
R�코�ȴ��a���i4��I+d�Z�$�O���z�۰X�Y��-���D
5�Ha򨨴�u�K����?Ұ�����r������1�	�z��2\���iј/d�#Y?+?���!+q���f�˯����:ZE�u�W�����%O�[#;�u"x�Qf�@��@W*:�ۘ�����@�Q�`�B+�p>���&ڰ�s�ܴ��d&�]v�%|��9�/P�%�mkJ�o����ݡ���M��G�g I^895���]rE��s��9Q��8R����)a�KɬI��jɀ$V߶ڙ����z����*�9*d�BQ�K�i�������WD��hp{T�8k��%��r�|�\��u��<��q>����8m�_��,g��i<L�v@�9��k�;|/-5�4q	�Ʃ�W ��9iMe��8��H�n�¨zW�m/�_g�vҦ r:����5�$�U&����TQ<7�G~	]��?�l�J9������]����~B�Sgܰ��_h��8�
I�B�Aw'��� �o`��?gȤ�^�����1$���a�� �jDB ��o�/;@>�� L}�|�Ӿ���:Ջ��b2LDUA����C��e��=g>g�aj�,٨^��oR~q�P�9�P�Q�o���B��W���Xp�To����`۶Hۀ�rl�<��9�j��P�" 4}ހ�pM���a���b��w8ڏ����a��bt�˿>\����e�ۙ��y;�<�:�o8}d)��r�􈖟�.d��8���NjU�a�4��4.b�>��r�V���2cF�>O	Y-�%h�����s��jx�E��d���Gٟ��d`�	��2� fjG;���L����$�����p8 .���U˨n�2�Qf��-�o-ʿ�|]�Ӑ ��J�;T[���{�T�[�ߖ,�ly9��r��*��Lf(��i�K�S�Vp��E��yK�3rsT]ȩ9Tsn#����ޤ@]j^��{3��a��W]�P�u1�jd'�6�e���" v��,��B +�GW�z���E��4w@��5*�F����nzT|�^��~:9:��d�'��I���c�3G﨑�B�>AD��G�Kԡc���s�c�}�~�[!m)]I�Ȅ���C�M>r�'!gcJsvق'�ޡY����?q3�b�gMA�_Ɠ,~=���5�S��>��=&�+$zpuNHD�	�
�̾�ՠ��U.F0��ֳ�8Â�ש_�	A�s�ד���8��&jc�c]���Ś��q!I%��ʵ�~�K�'o�O޿I���mC�v����I�2}G0��}�0������	�ڬv8E$� �c�c�s/���USo���M��o�>���l����hAj;�M��~�M/`=!l-�ܚn�����׊a���І�Kp��#��t<K"49wi�}�q�r�6���؞�p(�D'��q���p���ͱ�sD�t�g5�\�B������6�dr��{�!��569��g�Ob͵d��uC��@����%"�8ABtq�6]��ij�:N�r�,����z�� ��ĐY
b%�������O`���J��PzO��K�.i�ꝣ�L[QMߒd������%=�ﶽH�-��jö�w�JĂÁZ�E$�#�b��է �»�'�4����{,��y������~yt��ςDxQ�����i����&�m�W �*%��%�sztD����e�p-[�!���R�~o���k�P8���3��ע�S��"˝Q'׼���F4��ӃݬU��� �o	���XT�$��{R	�
"T���Յ�j4����?�5'�l���s8(O�x� iBL�
��-J�]��0Wѭ���Pyo� ��:p1S����mq�TL=���Cq�2�fd�ɱs�ҨQ��> ��͉�D�Ʌs����H��,��^U�AM�T�Ji�,��/�=�����Y	�n	�K��V���f`9u��l�������B#��7t��~�vp,��n�qKG��w��rr� *+�׻�
Ä�^"�,LH=X�3��@"������+u��-	�^��#����A<��ݻ#	�D���Is��2;´�~��{l����r`��U��cG��`�)������nRӊ�Ic�&'vg? .���	֨0�a��L������;�p���
���3��WR�����6��$u�7`�����G��t@�.#�*��P�l��@����.��C�̀�rr��[-W&�^u��1�='��戌r�w�O_ʵ��m�'��9��KmI������7�xwd,��!�kB��hS���DX��zI�;u��TR����kA�?lܕ�N��XFRp{��f'�,�V�̗�z�@��poK��Munyak����v��/`V)�Z�u� ��Y7SJhYҘ3KS�����8ܿ���8�4K?��� t!��O�C:�;�"���u����
68B�2���LB�{��u};�E}�)ܵ�e���/$w�ʬt�-���%
�( �˜�u=s���1�����y�}6�d�Yh#e����&��V'��j�"Q��OE�V���S���Jdn�+4<G��	/ɖ��s�5�[y����Ynf�V���?�[k7�F�N�,�66�?o8�H	��(�0��T��[U�<���i�j>�XP�~�{J�gW7N۶]��@��l'�\\�"���AF�	w�}��,Aj}/��~���Icȋ;���a��Ϭ{^|��-`1��w�<�|Q�v=d���h=9`���o��D���߾�쳞VOs�:~e�	=�BRǉG�)�V��n�Q3ˢp>j1�Dc=�[�y���
�<�a�o�P��VC�h��n��מ0Eke�N��k(��tC/p��bי���,/�j#*�T�'��Aь�~�%�w���9�ة�|<�؟���$^~`K|9��sP�'ױm<���Q(��c]¨^����~c`��3��a˂%�iZ��.���X�x��dw���i�<�������\��(Z8<�����|��������
�\:}Yw0�)S�.�G�/+DscN�[6�4\l�Vw��- g�"[�=�d�.����M�}cݠ}�돼}��@����(1��?�!����;�V�m�9�@�[�����a�\)�z�#�0���&�����W~Tib.��ȜM.�\���U�F!�5�K�;n�_P"4���̤����G2!�mf��hz��F���jm�Y�s�Ki��I\��6$�-4����a��>�l{�iw>���ZC��xr�6i|�c@��A�C�<2-K&�A�������@7>��kGÌ��S����\m@���ޱ��2ޤ!�d�W���|�q!%�N���s�|���1_�>���|����%u<ѻ&uZ�RFVJ7{��AB��t���ב��� ���I���㔼^���X��6����ADBx�Տt#@8�F(��*����JBz$/��hPF�7B'��D��8]Ì���9Q���#�&�x��g��k)����	���3��r"��L���i7��,��8T�c�ռ��X���LxA����ʸ����W$�~����k��Ib��\ě�XJOo�Z��$u�2*_�������]�=)_���e��X��~
L���S�S
�Ra����tZK�pygm]_2!J��c�BZc��K�G��L>o�f�m�畱��M��v��D�.2s�b� �x�ȵ��T��c��]kR�x�
{&�y�ob�ӓ[H�2�wE&X�Ϸ����UI���4݁�D�e��`�_b��c���*�g4��$��h86�H�+)�o�0�c_ 2��C5R�=£���$��|��2<��W9[���	�'�H��ռ&��ՙ��f&j�$#�ǜL+f�bGXUt2��y3����^�8��8F9�_������٤��&l"a�6�M�/�͖d�ޡ��%o�/\�W�D�������!�jE�3�����#���A߽�wd������IG�WF��eSR�g�R��9(*?��&nA�kƓ�1���9c$ݮv0_��N��Y!�
�4F1��o�$۶
6���-�1��� ��=���w�r���J|��_���� ,�-q5�9!m��P���kԤ����f�9�P]ce��/8v h,��!a����P��tׁݑF�H�5��0�50�qgC��q%&��"�I�����Sb��Dl�}2��e�y�Z�����K���.q�Cq�p8(F9_$�d���)�<��t��0�SK����L�\y�.B��q���X�V|�E
��JQ�,q�u	&x�|� +Q���ĭ��������${����fG)�;=�f��^��}��+Թ<1]�`���<c����/7�3
��+�:5"��'�a�#�1YޫX���Ҹ�m�|�)��_Rg�:�����i��6�C�4T,D������o�~kC�j2���$��ݿ���Y�Z�=��p%;��vr>�yĐ	Ԏ`�XQ,j.�Ѝ
K���*<�o�Z���q�n�����b����i�'�h#)�]�~(Z���=�iltVRv4�}�G1��@��ÜAJ��"�J�ۊdK���;b(�g'hb��fn2C�U���u��Ƕo3�[�FY�#s�S�t�e'm(G 4�mZ�Z����� ��~��)���X	F@ĺ�N�:�4��Un��)�&��ȝ�Z9�B,^�~ug�1qD�}�z'��{|�?e����Ѐމw� 2��DW>՞O��M�Ή<v�|'��������H&E>���P{��&	z�����Q!���J�����x0��q��%�o��yC`���z���
�#MZ��H�bZ7��4�v�+6;����B�I��&4e$��4n�t"��.Û�LX�p�J��L���0��r��S����T�w�/�iZM����J�t�����6ڎ6N�lU�����U�VEW�=0���������~Z�2�z���F�X�O��m��F6��M��+ ��Lpc�}=P�#(��'_6,/r
������܀�0WgP�C?�ɹ]��8:j��	�h?V[A�l`q�9�!������1:��g*#G��<Ԡ�:o�
+��ō�[�OF�������~�-*�}a��GcB��v�v����b���ᏝAb�%c�2'X�\�eR~VK��9P�K�����|��q��,u8�}�2��Z��;O�t���g��g����]�L7�/+�O寂���P���u��'����tD�C��RS�}J)2�����b%p�#�m�5��$�F(+v)@�݊1��f9�����CFUh��ت�A����@�z+����`�$��y�ߝ�˞��'f��f_�Ѵ�?����/�����->��]��׬�vЮ'�G�W ��f���hq�?��_�j(��\C9�i� �r��=M�YH��mK{ت��-�_z\�kOI٥4����K`O�Ll�֥�Z?�����_�"b�l��Fy�a�Z%۸8	C!���S���c�}zu����^����aZ(�ĺH�۔�Z��v-R�?gA����K[��Y�����u�~T�K	���&�(A�:�Q9����L���� h΋��Z�g�J��B��JV���a��1>%�Rd�G�@����+9��o�����UY���W��4�0nc���:X�A�*yj�5�4߅�t��>���P��������9�Q�	���_noO�A@�:�� B eR�0F��?"�L��dkeJC����%��'���J�  g&4Z��#J���M��ZH�ipDM:$�L�%�
�V�n0;��}����
 UV)�ڔ�'�� �����P��Jw=0�m�>����HYӓ
7%ez�Wn&����a(�!�����]#���uX# �fG;q�h��J�ϪMG��ڊb�z�!�=f,)��1����c���ֿ�,�_��������=跅N��R�C�� .c�������>�"/����`h�a4��J�BPh�@9�I�G�Bk���6Ǻ�TӬ�ƪ���K;̿+��^��h/^?�8D�̀m����4��;�Yl�XJ�SO�wu��ۣ�ɖ����,j;�ժ�-�ii��I{��.��>@�`a��pJ�.���t�;{�%̦���.,J�9�䥂�	�}z�di���T�?ڔpK��Ð�t#"��mQ����r֋^�����kB�Q)my��p`>���rKv�H��m�hlk�t'`Ć�<��`�J����a�_�91��Z5���C�cH�֒:��D��~NOB��o��?ê#(���Hp�S����`-�5���L/�H�3%�N<Oµ�}�~�b�ݭ��}�i3��	�M��6�/>	|9��蠰ݘ���2�SI�*�Lju^��p�&�&��!Y47���H��Kz���rCa�"�!/}=!b��)�ϧ����}��ܯ�#��j����>��X$�6�]E�\c�͂�?}�4��̺N)�I�eO�.���p���w�;�Qe]}wɾ5��ac�����	�`(RI�p	���Ql��1L��fQ<���!�Pr<��3j��~�?RV51�bx��x:[����N�$ES��c�=�M6[0?�#�6�z+-� ����<4+�%b���ȸ�L���Q�y����>���QG��(�I���]��\p��2`�"��fc<ӵ��UA94Ǚ)���+ ��u���F�#1,�/G�}��9��,�#:�4�ԛ����̜9�:U �sPritdUK�7~J��G �w��&�#+�Y_�xAZ0'T��.�됃1�(~$�W�/�@iÎ����G����\��M���0��'������)F���[p�r1�����~F��*�(�&�2�!�_a�_?�<�P}��J�6�T����>�eP`'�`R�Vf*e\)�(�ժ��`��M����<澐ޝ�?qw/,8�3@�H�n���wR��i����4CSAv!�ָ���R�_`���2�tI5�u>+�̯e�dm�<�)���K�k繠���P�\N��כ#�{�+:e~C��<=���=��k'�h|�ᜂˑs�?�חVq��r7ږ�z�9^c))�,+�:�aoyz[?���4��Ct��\�tSۑO����蟔Zc��l*�h
8�;�d*���H(7�S��M���W�θ~���}	����(� R?��y�/J�Tto�2�D�숂(O�EhQ״	:?u�-&Г�$�L��f�}i�P���r�K��` �x�7IҒH��5>qF��h�:�j�^MW� ^0��_a�?��O��/d���?����V�W��LIJ!Dp4�'y����$Nc�7=(\da��e�d��_/��X�yX�Pp�D^S�p&gÜ�_p�����?mk]�ɼ��S֓>,��C|���
2����r�����N�n�y�',q���� wK�Ѧ�M`�:��]�$cb゘R����R�go/��2Yyf�������?Ȱ�n���.0A�Y4uX���L�)BS����B{����k3�N@'�/u~���j¢|�<��2���W�
au��/�6/]�ٽ�ThLo]	e�R\�\�_�8+/+o�������էN�Q�|@��o�#��m�"��]C��'y2��W�i:W�{D6rZ��4����Y����g�S�� ��)C��s׀�x^Vc�ՠf�o���t`�:M�@��no����;��-�rW�ŗ(���D�U���;@t�A��ɮ��BoP�X�y(���+�(fwo�Z�}�N�ړ�4�1.���Ch��Cٳf�s�q*-��2p���0�7�������@�rk<Sf�WE�W hDDl��;X�.�{����C���v�am�C�����i%=_A �Y=,�<�hSv��SG�V�����O�0C<�B�����y�2<��������Ֆfr%�S���M���g"��@Գ��R�U�A��A4>_�� �A�WMzRY��uZO/"�w�.�_>дˡ�HS�>�
��~t�C}XI[�E(���zx�`i��+�~'���[t�Y�d%K�JҌ#˘�C��^-���6J�- �jq��3�8,��-%r}{H���)�Lh�gK���q�@L3-R3�o Q���У\3,�v���)����EI]ئ9�&�6�dBI�mr+&����}��I��J2��%�Q�$n	�-P/�5�@NWč1�x
3����Y
i݉M�u �)�AU�uc�l�a_u~��O�0��2̆�o̊̀��K~�����N�ѹ���y�0	3dq� Ì;g�A=Խ��N��T�⼂��P�W��{�D�ܚ<}zu�����n��1A�����/D��~��~1D�X�e$�E��/��a2*ކM8:��}�k`�x��c��~9��+�XɳV��i+|hm30��ݸM5���e�;�P�bKR	P�_�a
�A�"t�-+������{b��>�R���wl�H�7
Q@sjا�^,��f:[��љ�|j�N-R6�F�#n̚��C�����ҳr�c���(L��BK*6Q����������_>�~����|����g����EK(�p��O;��F>����ح��N;�LQ�N{]9�:j���2Km:	�Ǡ_�{�KR�ι�7�ĸUV%�'�3s�Qx���(��n�å��n�$���W�qH��^�̀G�=OC'mP�Z��x0�<-�x�B��R���軰�R�`���/^)wϮ�($���Iv�����e�V2N�h}���;N��}�ġpo��%�2��V��c�s�m��F��؆�g[mq����_�rN�n�K���MmDya��e]�B��4Iy}]M^l�)шK�S\㎞��-�����2�!�
�<�#)
ÉG+�.i�睊�9]F����g���0׉,������?Ү�WF%&���{W"�vR���
��E���5���~lL��U<��nv�Lm�� �&/���A�~���|�ד���a�8i&z��7����j4CJ&"�S�ļs��X5�\�s���9~u����0,� �����*���$i%�d�߬&�B���Q8�c�Wg�ȸ�i�������c�)���$0���y�ӧ�k�B�9�{[}Y�>���rI�u5×nA���uM��s�Ik�6�m��@�*0�(�_����.���]cfѷ��N�I�a�7t��y��.*�NvF�D�I'�}��?L�� UdxQ(�<�O0=�$���0=%�lDT+�B ʅ��޷�4s��x&0R݅��Π����Y�dx�[E����I�&t�X��S�����zC�?�%�~���L4�O+32UE���tX|�(��ݮ���]?�D\���+�l�e�P���x�-Ds��<�s����4��G���N(����ؚM�;�uF�Ô^lԇ��J�g�-x�\����BNx����Pݿs^¸;�ߖ��O�d��
���.�y�+�H�]UEO�}��f���BTZ���iޥ0���,�\�#�_��b�v�P�|��i�P~�BP�c<��桍�Ji�~A���}�����v��h��~,��~'y�E�ԈG[V�����{�I�ӱ7�ҩmS{,��s�%饁�t�QO�/�S_�����\�? ���hm
Hj:!${c�]!<PO�����Y�Q�`΃0>������5�J�AT�Uf�g�<Z��ޖ_?�\�=�A�@޾!'�jN��vq~:ф�3�AS3�Q�-�c�=[%)����y�N������2�g�/wbl�]�w��RC ��؁D�H���Ϟ1#-T�E�y�'��!���&�$�������ɔT�T����yC+:S�b2��a�'�Q�Z�nRT:��ꅩ�)���Vb��`�q+8�.N�6l0����;$ė�Q2��r�H;���~"����#B䤽$J�Q��i�nAYzYJ�ሓ'A�^�t���49)� �?-<6�D�=��E��%��O�Y���
��v�&�TϤ�A�O4f*��a��a�mս@3�Ar%�G@�r�N�}8��
�կU,��u��d\�p�˿r�k�movo�W�
��������o.ڻ,�t��fH}��W�n�H��؆�Fѻ�O�ޟ��t9���:�[�_h�:�F�ŕ�0_�U�⪝lCkJ���!�k3_�~0��m9rx�B}9[DA��R<7�a�˳]��O� ���������+"r�`Z�����X
^�	�ԛ�ٱ�}��#�d�J��-�jPC@��C�7����މ��_��n(��S��	4�dP;v�Go��N�ũ��i/��x\�f��|�E�Ǧ�.ϼ^����Z���:Y�M&��q�Z����"w?DT6&,�?*8��(G|z*[�e�. ,�l�Lm`3fU�P�We"�U�>W~��I�ג������N�ȇ	E|~���<��~���:��:9�<��&���c��r������t�����OL�h�  �LY�bX�V��V����'�������s��!߰-��7�HL�l�D߆�x�|���gt�Z\E73���6~�z�QS�%�� t�"�r3F�vN��IL.�c�wU硘eH"}R8�o!�����glj&�b����`����?Za���*{d��m]�l�S�P4!�l� fl�O��?�xi������7����?}|�.�B�/�8�NQ7`#�\�S������;`�m�k���.�9s@L�$�zr~���i"HM���H4��`�A�U*^�b��5sl��qK��+�2��)��>[F��ް7�	>�6ѿ�5��lML��}3��"V��oҰ��PU�o���<��FLXI�ѡ��A-���6ui��oO�/���5Z���K��hFs��~]YT�w#�g�����%���؈
g��]4�~�-u����X�B֌.9�b?IE�b�P	��G�YzA�H�Y09�\eR���Ȼ�Q�d���et��q��ݚ��_EbQp/�6�IA��	��|��T��n�g�ɚ-x+O��s�FȒ#�>��=��q�AA�9�߹`���"�P�<e�2�7�	��t*Q��C*dB�4ш����4O�8�RY�[�?v��aZ���>�v�h�9�*�.���f/=*�����D֚jvk.+����a����`���t����}��|B�>�e?�h�=��%=%-�e�t�v}=g�c������&vr)C��WȀ�6�F�$�<:'|V^߿!`�Z�����N8��ի48�
'Zjw�#Δ�2����v�k|��HcF&�+�1H]�q���O�ط��q^���� �mJ�4&�������-�O�Ȝ��ʅ��2h�9�\���^8���0f
���d������S��DX���S�D��o8e���p�5�%w������>��B|�����%KYhm�?�)��B�p��n'��q���uU�n=#����EhC���D�(��u�k�%�*�cy�`$Ҕx�m��ˤ���u�� �<+�T�9#��n�fS���ޞ-�]h���]B�%N3Y@-sa��3��*�q� }��7K���|c�����}9����
����>}� fW�f��c��i�#����|������ݎ^{ë���K
�5��T��[M��PT1o�J��>#<,��؎���� �~��go�<B
rzU�?��-�q������>j��+�3Z���x�L�T�Y&�i̌i���4�gĲ^��������V��6;���O�^=f���R��f'ϡ��S�v�\�>��M���<V�jU��?ޒ;�uj�?.r������\r{��\��	D����4�_�ܤ���1��cK���\��^��*:��uW=���Ay�S�)oL��d���* +i��d��f��3�8
�W�F����{*y�z��[��-�����׎Ip�9Uu����X&�n1�$y�z2E�B�:pƚ�0Ŋ��5���zR�LSX*,��d���F��!'Yh6��C�eL�f�k�"��8�[�ĵ�>��������S^�m�t(j,)qh�~
�j��E!�f�-u|_�y�$�utǧK^��[��r�)�����z�sX��K9�m�gqUl���*l�-���e� c�<(������ıI�~� 9�D�I����
��Hgo��3�*�5yO�.�D�K�����_b�:ف�;!+��[Ch�3��{�塚DM�,���-�1{���'=�� �@s$�_Y����I�0pK
F��� `Q\�j�>�o���y�e�����I�m��]�l�:�����lL�m��^�����Ic��z혱�6�)�Q��.�-��*w��뽪|�kRA �1yT13:���iQ�T�%m�r�*`��k�}�(a:�Z��pQL.����^qO"�<H,�v���-�����.셠�T�A[7�&;����c��7��[|)3{��D]�Sd�ja�8i�g;��d�I���D��(�j�n-���C%���9�&Ā,�=�~�L9.7+]w.�1UБ ~�`���唓�{����!�� �`�����0n�G����Ɏ��DMOQ����#0��c����"���/�=�j��J�\|�J9P)����q�ҳ�\*��k�rI�R���	Gʀ�G���ύ���*;��
��%���e��t�a��\,{z|�ʩ�������~�����O�� ��Б󯶒N�iϣ��ؾW�Qx<ւ���qL:l0 l��w�K����'N�1���A�T���@*�$x\)�>j95���a1�wO�Q�z!�ֶ9b22��x6��g8r��S��Dzh��Nwf8��g�XK�oL�]��\~����0k��j�G��-zDy�J#�bu-ˣ�W���(x�r(�^ ��T�3�*�gO$�9~��`�> �DŪ���M��Q��!;�9Uw�o��H�C��ob��K]n�\�����m��}�|�*���9��HF왜.���$��H�'n���;�����%#��=e��'�:�Q���,Q̗���&J
g9���7�7Go����b����Z�r:8>���L̪��u�����m�}O�d�>�)I�K!��'(&a�1[ي�"Hj��k�����IԔ[�ux��Czg�|�	�S�����c��"��Ԓ2��O�]�h�5 ����fU�+[����V�3��Db
MN�Ę/�C���ڇ��t��)���j"���y���~���} ~Y;w�kX��Tg�!�<F�w΅y�k��<�����ٔ�.) �@^�C](>T X��K�-qA��3`[X\e%dt�o���r����;���	����e��\�1	�X=���p��?��pw9��;z��N��<������mDg�������@�:69��ux�j_��P����h�XMy�d�*P�c��;�c�<��߱#��֒�k���a�9�B�oϤcδ�|�V�,n�S��fYY>M)��u��"i�|C�heQ��B�N���L@iמ �O�����c��Ԗ��Ӎ�-���rzVm��n5M�v]��	���tW5���ōS��R�ɒC�~1gG�P��~�+p�t�l<�"�i���դ;Q���^�V��(d0��s��Y^����,�w��ϝ:��`�����nBu�2Bzތ�3���:_9��*J�p��$!H	B��E��km����Vb��o�V�ոn�V\�H�}��Rz�d1|�<�c�:Ý�2o3��99��Bz��j 
r��O�U���y~���Z�d�J�lǠ�֪���_��
#LT1��)�>W�b��8�m�s�50:�FQT��������w�P���s����I*g5l!c*�
U��[8��i,&,��w���� ֦��kͲ9f�.J��>!�ˣ��U��PC�ߖ���'��������&�g2�E�8e� �:.���T��m��Fw��"�z���������E ���^��$�kj�v	Z6�-���(hV�^����vz�5�pDy�4�O0w��q�����`k��1e�/���W=t;��o��Y�U�b�B�{�dWO�c�p�Т�΅��pKmbR�ּ
�\���������xv����Y�g�ߤ��d&�}l���m����8��o���U�����J���k��>�2������"�áen� �����ʄ*�sl݌5m���ZҴb�M?�����X�������rwffn�f�PG��M�����(�	F*g
�N�lG�&S`\�F��c�d� 8��֢j{[�6����Ky��xK�'f�&��f*�K�`�
�U��kR�[�{~Ϙ���� ݰ��c*�ޞ��R>��,1I�_�;k����8�Ȋ���ݤC�X\N�J �O|�.���#X9�#�?_��[��{v��㨩�i��8Jl(f�1�2�����A����G�b�,J�����K�Av�wG�7h��vl�2OS��2<�?Mػ���6/�q�i>y6d�"�]����RR���(��~^@r�^.i�����#����+��J�������/��^���#�vTb�*�!Y��z*��������D118u��S������yY�	��@;;z�8-X��Y(#=3;Q�Yf_,�w�rL�m� ��겓����N�V`�~�P�Ő7UVJ��},\�JRwD��0�/�x	����%�(�Ǔ�z�p���~,�#/���h��V/��
V�E���a��d����r B����&˙K�Y8OU`zD{_*�0�ua1�,й��oV�:9Xe��B�]�0�]�r���Vcx��o�" �w���3L_�=�2C�����/��7�|Փ_�N�����{��L]u�]��O'�^Z�}f�B�(f5[c^?[���"� 1p{is�p�����d>(�����䅩b���щ��9vJr�GV(�=�Lw�E�z`�j N<a��JY8����{@9#;	d���Y�Ų#C�sz~��Ȣ���뜸�L�>E]yٺ�n�̡�i�� l����$x��aV��g���~N=J��4G��E7��x����H�X�:&���j)Q�`�+v%��y�������]�\�rG?%I� {��%M��";����Ǫ��j�qӳ�T����˂���A.�!ޯ(`b�7��p�E�9[���Z���l��:���ſ��hOLFDK���4O�
�e%��ﻣ�#E�6���Ar�=%y�ݶl@��frV�Z|��S;VOχ^]���ʃ�
IhFr�kB΄��̺;�� "Q[�`�-?k �}��f�`*������1�`X\mv�1���F®	�3��n��鬺lD}��L_|D��HR���fM}��jO�h�0ҧ.<��t5�f�D+"��if��ϩ�qp4v�wl��<n|I��7��x�Mc����g$���J�ՑY�M鐪֯ ��1�]���������}���o\��)r{&�	�]�lZ���G<��-����QxbS/�2�@���c%aάE�]���́��Q1��'f��OiH7����ps�<L����}�}�O��c�/J���`��\����
�yH�Ŋ��m��Pb,|�M��ҽN�Wk�_%�g]�im�87����f�m�ouԸ��Q�=NT�.�i�j�	jЪm:��� ���3a"���K�O%�yO�_ɏ��~N�q3I��ýk�ҏf�r�p.L^/�e�aEE2Mڅ\���{70��'�A=�x+��.:�Q_������l�=v?�~?��� /�K�M_���׹%-�|�Pl)�4��Bᵾ��Ҳ���ݮ��L�{��Hg��< y`1���7h�� -wa�����yE� ߺ�����	�Riw�#jl�2�xޑ�>����=�Uh`�����<j����87�����y��2Pk��j
�D�1���֍j��[E"�W��ݛ�z[�nA5����,�x3���o;����B�-P�W ��0�+��.N�f��9c
}Ĺ���s)և?+W�0��"��J!�+a+W꧉WU����9��.��Z ����"�{@6 $D�:(�,U$��ާ4�iA�#_�	( ��`"��;�d���wt#K�(��x�2�f%�P|�@���5��NZ��9x"�4��vf�XB�Xҕ	)�$�7�^�f72]��)�+�**�)�DM���3Ǻa1�z�)�j�o)�ˈ�8_���L�=��Lw5S��:w�uir�
nMm���������KѽR��q��u2�0�6-��cJ�K=v��`�8"�9����p|�gjL1P�j���m�%���8lD|�x����j�sr3x���20!�y�a��&�/��Սs�����[X�w^9v��_C�}��x\k��Wr�����҄T���x�H!䉠^Ay���/���#��~�l|�t�X�T���ռ\�Y���9Y�^gz�6�9F|�r��q�j��1�PY�Q4�]Um��{��������&�	Ye(��H16���;往p�'߅�UM�?F��Ŝ���YV���+�k�B� 6pƾs�
�?[�ctl��Q���7`{&���$	wT��|9�;@u�]��)�Y���uۋ���Kh�q䤡����f����˾���d#,Sk�Br���΃h�vzҼ��FL�/�XA�|+����|w�H�z*p�c"���3�F��3���$���R�9�=m�?�0Ϻ�����Ƥ�|����H�7N���t���^�Xjupл�G�����e[;��LU��۲EP�����R� ���ަ�[��t���Y;�$�&�����&��i� ����f�õB�&S{��p$H�S*�5/gjs�-B<����U="�<�l�Uv��|K��Z!Pe��� t�oD��U�!��N���Ppm���I������d3f�=V�ܹ7�aU{�>�ն�G4]��K '���vɥ� ]I��!h7�bɲ�M��P���2�UC;�n'JWد�dH���	�0��?�(+X�E�I��%f�C�p�����$�؃Y�)w<[��*����ݓ_�ی���W�����a�3���'Pe�ȗ�[C���:�'��c���Ԋ�i#h9<1Z���S���@�;Cg�g���:d�C���`˔7��b��HH���z�bc���Z��;�b�sin�d�V`	˘Ǵoz��PĺЩ�pzZϪ��-y�v�W�K>	dN����O�N�c����B@!~�ڙ���tTf��@����Sp\׭	� 	qLw��3*�3��}��SO��;�WŰ��+�ȈD�J/�"�$Z=�i�.�@�� �w�}o�f�J<���)��0}�~���3��0�x>D���ge��s�v���p���p�@�!V�?ɉ ���s�<)�	V�"	��MƆpI��l�k�K��%�t��@�^��htiP>Y	8��'�9e�-�S�	z�ލ��.i�p��:z��ƥ��� b�/C���ď�E��E���!��UhH`Q3ڹĎ�o�
�L���I�2�@V�tX��f}W�۽�ts�Ӧ��$�ڹ4"l�`�R������y��$�]f�Ϳ7��)���m^��a�yp������ �A��XA��jS$�e"4�N�
,s]��kX�<��w������i��QS�w�f����r@#��9M�>d2�>�G~�p	`?3�3��$[��[Jg����Qc�O"**׿��W0��$�CZ���_��4��o	�4���r��m�����+c��a她F�ג�d�d����4�Q0I�1:�Ƽ�I�X�e�"5��@*�F.ڜ�1ov(��9s��D-s����+ vs��o�t�j�A���a���R5�+�
����j]dO"�V�1d`�xT��09x��������K�2���F��=o?}�JW�;��pL�Q�m�)�َU���J�[���c|
6��\��CΞ2���eÚ���L�g ��8������1��)G��,�������ކ�qE�<�[FZ��m�4��k�bb,wƉڙ�QF4�!������~,�?N�`�0C���\���/�g��r���(���h�e�9�۱ˁ�t���tǨn��w�U��i���c�ƚ*eW���69_v�Fi닶U��1���`�>8_�%��1���\�Z�%���RB�g:a�߽+x�ٶ��F�A��Qq��L粄�C/�r�� glt����X�
�?��5yEt?�:~W�~�������肄e�?2&����ZY���a0�O]���f��kݚ���WhC�B	��?H�H���b��� �Ց@iře�H7B��a����0��o�8�RG���$�լ/<[R���C�̕���v:>E�m�x<���m��N����w㎫�/���U�"FR�kDA�o�S�J����>��VX��	��G�M�U��9`�^	m����V�hI"sM�=̄��j���p��,b���uN:�:Jq"�{|�E�Yr��m��-�$AF0s�	�<��Ȼ]�g�prd�%U;���R�������ǅt9N�R������f�=�^�C��}��~�k�������P����q�$�L�V� w�=��c�c�K3����p�$����@+�G����֌�qg����2����z@`���������X��8�<�v!�b��v��i��w15i6.IlkF M��-#u$\<��_��8����a���c����u[�ٙm�>9�[cA�8��|l�r'�S��s���	6��gҘ�v}��͓�fF����I�����U�@�f�b_k��,�y&XcLz�jnC����T���8	���x5� �>�Th�B��	3�ۅ��A��M~	��?�v�0±:�}���b[n}�T�.��:�x��N�J�ւՓ��Bdxց���W�-J��Ɛ{bd*ym`��Sq˿���]��B���;��Y:X�j�F�xc{�3���>����Q´�%�.�7�XJȬ�@�ʍ�f�;���K�D(��s���;� #�T�:�����6��1��0D������2��k��H̤�2Ku��<B: &?R[g��l��u.�ĪO�8�@]���������{Y��,
���]�!� մ�j���{b�}	"ΖFl�"�θ�`���1��mA����8�F�Ҫ9Wq1�B����'�z��M%���ጟ�=.���5���nN7���{�B�7˒̏�����O����{/J�ޓߥ΢CfD�L�C�c��wKF�݊�y��P\���,�8������P���N�y�8���׏Z���%Bӏ�YN07(��f���������ԙx3�C�D���{1 {�=:�D\9�^����W�	���A%������2}�?�v��XM��oڥ>�B��!�Oow���ˆRS���Wh�3�b��61nԮW�a寛���`�D���)��\A�i�	A�^�k��*`;Q+�0��ȟbbea�/����	���-�?���=�����k�U�m\�o�+��N,h"v��,���N�aSC�43��/OV�p�(����:�.�
��?�7d4�ˌ��b�}��	�ϱt�s�$.f�&x� ���jhν*G�H��|�H>
�7����&��<	:��/��S�Oo�A|uq��-.}7�6L�	�S!�7gXWdL 6�+�A�	( Xz�D>��s��&妨����7U'�=���x��hjG@bG�j��j��g{��	1��8���1��5L��C!z�l �,J�&Dz���`�u$���:"����l�Z9��+���\��@1�2��o��~o���l�ǟ�Nw�U����|m���jG%A�}��1&���_jp�nrQ*�m��E��X���W����)����w�gҐɕN��>�ӕ�z��#��7]4D����0ĬG�H��ުF�7�CI�g��j;ׄV��bę���BZ�a�DZ������+
��F
�M��q��m<=&渜�4{�B�P_"Gk/�>�j��8�?�[_ǝ��GN6�
+�f3�1���D����^���S�+0u���~�Kp���^�F�F͌��W��x�Bߵ�<��s�`�~&	b���g[v�;�� 
���k�-I�W�X��^�֌�1ȫ����h2�,�͗��ܿpP������}n\��c�eZ�$��I�3Ǌ�Obs�Y^�<���MC�ipM��u|�)���A"1cB�\a�ڮ�(���0�Y�'y�|�������l�s�@	��6�qd�#Do����h�VZ�"�ӎS�����

2A�(���,�č#�ew#�d�d�
�Q7�m+	��;�`S���FWN�O7g�'�Ro/"Q[<YQ�v R� L�w���O�ԛ�T����^�PLI�͊&���OJ)֦PI�ْ')W�Y�i��w���� �������E�;u]:�1�9�V�0�'��c2!��Oِ�Xo���'=}n��}�q�w�vi�����w�x���5@!����E�	����4���Ia�(��� ~S*�� sL�S*C�K��6���J���u_V�������٩��,�~��)a~?݉O�鮬�Grq��~����3#��B	�$l���.�N���@�J�Y�JMsh��?+&'�eS�&�cck�!�[���w�a�P��6p���)1�nVǉm��Wጕ9h:��x�*�-�v�J"3'�J<BWn��?�SyB&6"���
[�a:c��)��p�	@�?7U��Ϙ<K��3:��˗
�W1A�
��ҩj*Ȋ��E��Ҫa!t�C�)z��.���}@�O���4�uۢ8Q���g��A);>4kM;�aha�v��3��׮�`/R�2Ǿ-dL�x;�*w)���y}���z<%ͨT챬�7˭��ef���/gP뚬-�ۆ��P4�<� g�@@-c
+�,@�Bu<<�Ј�����6p����@��E~_�����u��#���s�������$�lk��dM_#��4�gKC��7�!��Yɭ6a� �	�I����+�'7u��bA��0כߩ�,�[V���Qg(+m8�����%9��v(�`V�ױ��Vُ�=k6s�ub��6�;R�،1Il��͒�ry��Ά
��e�D�J3�V�y�C�G�w\��M<&����h��`���l�*�I�~ǋ�)P��le!�R�����}�刖>7S�~#)_w[z�Bǩ*��i��B������d=��Y�8�G-��/��I�}ĥ�� �Q�v/��À?c��Y_Z�
�V��_X���S@p�]��&y��4u��Ol4~f����r�a�Zj�M��t�Nd_yL[���$ʙ�H�����k����*�|��H]r�=��.�?@��=@q��iVi����޿u������Z"`=٥�[o�w٨U������29$�������k2�'Z�?e�~_�}��֮ȣ��; 9j�W�8��R@Բ��$��T�e�ϲ�ʍȫ��e�
�P�R�����1�lɁl�D�g<�O�I�Bo 1������n3���z$�/�����Ű2�lLM
%��d�(wH�����g&����m��8�w�j0��hF>sOp�\� �B�0d�8�m_d7[vមas�)��-l-��0�;�-�K�ɤ����}��z�HE�����	�F����ȭa]c ��8Ѯӣ�īw�a��V���Kײ��#u�>n��v ҁ��X78t���a�+5����zm���Vo���w7��c��wk���/]�e�����_&�ɐ�����n�$���E������J�K PEM��Of����,�>�[B�sF���v�PN9�kx�{���*QJ���#y��	 ����J�O��۫�l��[�M���ydM����B���o)*��@Hf�ɳ�L2K���?� 7C�	���D�	�&`�`-nYː��E�?�v�?uw�}�՝�� vӇīϦ^��;ts%Ǧ�#9	S��8�`g�q��6�N%��"��s�w����� *�x���{��N�"e��KȽB�d,ޓ����M7��]�}&�$�ƿa/X�D��0&���z�+d���I6�;bi��*�O��� �eL���!S���afz����ߺ��|��#��;��XHI�gQ_�{�iVx{��}撎�[+	pkq��{<���Y�fZ[���^�R�ќ�--��Z�Zq��$L+�#
��~��4Uz��)�za�0�{H��
�����.ܥ7�O��59�$���ms� P�`L������+{t�\�e5���H�y���l��2I������ �6�0���V�j�OGu�R���E^�E�2 ����i�s)N�1��=ZG�ukKC�w������L�S���b�5�A�n�V�.�5���`'�C����޺�ܮU�U�ue����'R�A�(��iV� Dz��&�]��Ar@�\HthM'�a��b�R��'��ۡ�yW�T�Wa���J��[�h� ���m��MV���#�̪g�v0��h�'j�f��������Oz�#fxC˥:j�/}�%6l�
����J>��X�6?�b�s��N�����y�T��GW�Q�<<,YE��Q;!L̓���:ﺸ�?25H\W�37��Z�n�h��%�������Yl7 W�����o\�]����=!C>�n����c�f�?�Z:p����V܋������M��Ҟ�ڡ�-�lO����$r-��98'�Wf�E]뽖II��/����i��R�,�6e�������JRL�"ދ$�x7O@��_@�\U��ɯf94�MTa�t���Z/e"�hGџ.�����h���[����ӆ����d���@x�q
���r��3w�K�#����k�r�-��6���VZ���7_�Ύ��:ӣ<�V��4�DZ !��ش��%����q�c�!��fF7܅V%\���h܀<UJ����W�Y �]����<�ټ���G6N��R�*�*���X'�4y��m�"X�ϔ����m�Jw���g�6�������g�X|v,,耦�~�82�:�a�"�q���/���mi@�mRm��%GV͢u���*��2
�C߯�A�:*���%����[aF���^k�g:OοP�s���?P���Z���ݡ��r��t-;P�T*�<��5��~�{�2Sy�n6aE�1�Qa�Y%��U�w���Z�k�o���0[
,�}�V�	hgb�^�!�:B��@3�eayY5��LO� �7Ȫ�	� ���)�Ij8���M6�ճR�ʁ ~�ﱓ�SA�%�)��+�����$ɴ�ط�	<Vl �T"(Bi�--J=�W�C8��,z�!cb�b��5���J�@�"�!u�UT�y7��bJI�cA�g0��6��ޭ�.�@���n���nIN���L2�@��ڄQ��p�$(o�-�@;kˬ�E�#�L��������8�ܦ��ů�>cd�S�� vq�k��K��U�d�=�ǐ��$9N깑l���,��kIKI=O��`iE�1oM�nz%���F��\h*%	9�OCV��t�%���.X��&��i_��^��D45�r�� �ޏ�./���2�����ffSF:A�J#����&�.cG��`b)�~B���ġ<��u��j�N�km>Q�q�ݒ~�at3>�]H��/��C<(�ԃ}�R�*h���kʾ���i��W4A�i�-r�q��貮;��X�s�-{�'�VV�Ԟ�w|��� �U�ER���`��o"%<		����,#���Ў_���"�߫�.3����(���h�ąX\*�`^J��Y��Ф%�U(�)��.�t7����8���2nt�#�o�y��H��cB��������x1�S}���Hsl��rW��<L'��y�y�,���[�#M	wz�&p�S�O/*Gvz{X{p[��
�w�æ�9���1k��Y�[<�c�Q�S���3Zϱ4^�v�>*�H�Y�}xO�-ᒽ~0�'̸��+JZ� +R1�d�T>/Vo�n�<�ٜ(��]����?L@T�4&p2(�q%�}[�QZ3,�)�QsgR�>Tpf@<�
�H��C^��k���c�M.�PdZk�d0&.�[M"����R�b�g
��}oj�0�n�}G���`[�d�{��F�n�2���PE97���i�1�lY��'R�x�J���`Ge�h�]�nS�P@�m�͆*]:�ć˗2���0�˔t��q�����>��WB�v�[�y���>ň$�Ek4�=��5�U�U%B��9��gY�m�؂�R��\�i���va� 1�)/>{�p��
��:I`��bL�#��N��R��aøy:�C���hM��~�3v3_�����4�bm��c#� 4sx�P������*�u���䌙vhL�kB�E'i%�$%���(m��U2�j�P`��)ҺTn�a Fs*�<�����{��Ѥ�
+���7p�xC�^�G$E�������Һ�e/y��?T �� hp��}�G�,̏��������ܪ�����b��]_�(� �k`��L� �V����Ʌ�0A��n���=�O�J;f�᰷��t4���s�s���OI[���G��I]��d]
Ė	�N$���Nb._]d�+`��L\[nDa�Oկ����a�Ƙ��(:�^�V� R}�E {���Bw�����:MQ�����6�$�K�X�%n������$��;wT�<���&}�×Y
�w_�M�������DT����G�y`&6��~ōڻ�Q������WM7�6K�5^5� ���6}�3�,@�����&O+@/�y)�f�^��\���ᴇ��k< ��xr2�e^��n
4r+cܷ�4��)��j��#Ν����E��Q������L_�u�a�$�����h���[��H��)�Rd�bD�l���S8C��k��Pt:�@��z�鴚sr�x�Eb��Y��h:j��1c˝��Nh�7�M�� (�[Æ?.�!�g��v�/������Y��ST����ψYa��M<f�?�ͻ�����+�5�߼�z� ſ�ZK��4n��R���R�8g�{��6�=���x�g#��@X]#�]�5?��zB�k�1�^��6��9v�R���%�-��g�(�4"�KO��K��Q96�1�w�H9X�;�8�4~_f&^�
)�0��7����9!����KN"7b�4i��Go���K<؀�'ߢ�yq� c{С�Zz�J�JG�k�"�����$�UK+�M�'A�&'f=�E���)��l�~�eE���A�%��ay���_bU�{Uq��h�r�F	-����%��y����{����^�y*��.f�om�d�k�+�*�Y�0�� uO�L�<M��BK��I���7�!�?-�p�">
9���}�Y����<v�Oڊ�k�"�N�?�����U�S	W�������0�3�r���/���+`�1G�jh�D:�]���c~ßH;�6��p���ڃw=���>`͎�����(��ራ�����2�t g~����==�b�3��1�qyl�#6�~����s��$?�l�`H7O�"ф�IW�Î��	V���U�ኜ�Wpr���1L���������oLm�����1��Zd7���ſG����/
�1ǔ�ؔ���q:��
�����5%����D�~#�X�.�	͵��ȝY(,	p�:����)�����P�x���a�9����'�>�LN�13]Aw,��m�$��U��S2ȶ���L�؁Q��G̉�a�#:��-�6?Vj�!��!T��_o�#`.M>ٟ25i�Q���h?����/���K�y��8CYN�������W/�%z�|ԩ�H���[�2���Z{��k��H�%�o�pN�<��ߔ��{�Y#�S�����&1��`�ϱ6>���=�.��9h�q2�G" ֜�/�£�F�,C˟���emۣ.b���=O�,߽}����n�vz�(a�&�g8�$NA{c�f=�R���(�/H���.��L��x!wuz+)=��z�|�(M�a��-ւ�}��	�Q�r���"7�Ԃ���E������15&�Rr�KT|���A3���v�Iڌժ�(�yA�L��W��g��x�-S1Ѷ[w�+�! ��*1R���	̸h-�׮��ёi&;(=�V��<���R��N+�9W�E����A�j�K�Pw/�<��.��o~��3js�;>7��£��S͓֘���4�k�����>[Y��	�_e\$�yy��2!�9{$�w)��,�e�jU/,�t��2\���/����lh�+i�������2�Rǒ����V@��$��!�ǚ��R�W4&��ɬQu���r�	J;k�=�ƙ��x��!ܰ�Y��RW58�"��$TP[�_��p�����#���گ�B���b���&�x��������[S@w#����+?)��֛�O]�k�����V�����g5����M�	z�H�$p�����p"6>���%���ӡ�[>����h_>67j��pA���.uU�N����S�ې�v2l�|���k+{���a�N�"&tZ�w��?���.��2�w3h.�z�f�n�,���)�Wb�B�y!��RS&�{�J���H��rA6�y��N2-��/L�R�vΎ��9D�O�Oq�7O<*j���"z�pc�w&�s�ݕ��飒Q��P��:3J���ˊ>	d�&V97N�%e�F�e��.�H�
H�x����`#��*��TH���q�$v����m	�"!1|?	�ف���6�Mݸ��	S]���=\��c�}�2{ڢ�%�tH�t�R�����ZH[�����Q�8t�@��*E3���5��`Qv��?&�@�
*���܇�Tv�b8t�E���w8,�¾ D����e�0�C9��fd�����*����~�� T���|è���]�Q�h�[I��ax�6�
(��ABA��sA������}g��{v*&�vU�������2�H�q`�T���$�*�VS!f�?�J�0PYe���75t�r2N�D�̽�3���܎L�`Yn� �P+�c���&c@�m����^�#(�bP�+�,ˍ��b�����2��I��[s���	G��F��ޠ4��Yrj�V�����}�R�P�)	(��E�E]Y��GodҎ�p�8v���䩒����Gس&�I���
�`]��$�.�7�oӯ����l(5޺���X�{6Zp~����Q�LK�P���3��1���WyR�J�چuJ��r<�lH�U���GB��_,���Ȋ��)L*U��ӵ�)@3��`u�u�h��Ӿ���*�q�)sz�Ӣ���5D��/�XOd/N~�ϣ�ߗ��{�=��H�=��7�yR�̄���M�v�W���P�Vu��c6�-�¦k�n�`M�h�rdj��<��7�θ-� �-�d-�Emx���V�D�7�ꍩ\�{B�y����~n����:Ч���Ox�� �,�\�i�"�|*��lN�l� �_��)�"^�H�]�Yɨ�W���*s�������5qo��O��L�5I�I.Ҍ	*�| '!�{��O[����d�/f�^��Bq�9�Fc�t(��䩝/�ep�g[���w��ܸƚx���EY��/���HbShv,����0T�8fY�?w�}��Hˬ�1,;��,'|�/�&��%���@���c���(ei�N�K8B��?��В|2AݰR��d*Yw��x5���޹RW����/�xM��^����N%r(M �~n,�P�ǿ�T��lq7����Bǚ��^l^�����O,8�=w>�R���q芮N'j-��̝<P<6�F)�欷D���+�ԅ��I�v�3�
��<է�b�����D�x'I��y�/?�lMc�Ah�i_�@;�鈒i�5�6p����6�^=ژp��/	퐡�v˻�'�Ig�Kxii�D��.݂(c�:w8����¦y�pg;(��U���>Ƚ�jDk��V[��	(�R��2?�����yj�[�ÔZQf��M$PH��2n�{�y��M�ÿ́�jt���_���Z�H�-^�B�Azq@�2�_C�|k�TL���Muv����}{�M�H�� ~��Zk��EC���K( G��WT��;�<4�%�{ʏ�燳U�ً�-�P����Y�ے�/o9o̓��3��欚�m���]��]*V�����h��jB��r#��^��� �3B§�	cJ���A}��7X��tM��a��m��)1OЭ8k�bЄ�Kk�����:�#4��D$
����8F��;�����.b!�ϋ+�5438:cY��iڒD�7=U�5�ZS�W:S�"B��GN~^�kJ��J��g�tʖ&�n���LB�M_J$�1O�L>��K��롆f	�|�_E���؅r���W:�e �Ķ�/g��Pr� �vO�[�TL�f�4�ڴ.� lz��ٖ3L����*��"B��I�,- �;�C����-3Չx	a�{����?ϳ��Su��h��f!uMɥ^Y��*�i���S� ˓C�
�=�AB��=R��a��u�{�.���[���*���_k�R:d	6\J�4�Q�ew}��Q�w��Lg����K�Y�0Ⱦ�ÿەԡ&e��b��-���1���
�KSR�k�s�g_>s�B�c�PE�Y&]��w =��j�V�s��$�5���S��1�lYEm\�yr<^4��缿a��/���A�uRVTҒ�Yہe�='�3�ʌ�r�\wb�dH����x�%�B]p�qv{Ajl[�6����ѹCc~-%� ��%� ?߼��C"[�v[�Q�^r�,�I0z��&�?�|!G=�iJ���\@��t�$<)~9Z���1���i�Ő��`�t'�|E�C�/�M����8Z�
���b�V�ӵ�������"ȑ�`�]{�M<o֝ٽ�@�F�a$'�8h+�zD���@w��� �ض��s�p[�0��,����G��s�Z"rU�ӭA���r�[X�u�2
���f�˖y9���"	�.㛰�H̟����g2^^��(ԭk�x�M��[�U0o����D�`���ڰl�t*>F����Mu��jBo�����	f"��}=D|�����RG3����FLpv�������!�dB��}4��3/s&l�cL�Ȗ����G|v׬�h������rn.J��W'콽YG:���R�>�W�|cL�u�K_���dtv����p�7��M����PP�'�b�{�]�{�r_��4X�/�{�)"���𪋧P!\����7���3��v� ^��-�*�\RCa��Y��wуd�f�l���y�)"X4}C�4zL8�x�䐎�O�g�u�,Ȫ6�W�⽠WI�]E��֠�eJ���G;���fZ#�q2���^T}���� c��Ai�[�k	�^�F�0f��`�u��T��s�R�PI�
t	 �DI.3f���vgG�я�qq��3��" ?�)F�N/`v��|k��K�҇qһ�0����K��2!GBb�3�u�F�0\����hmvR�Ty�f����4ץ� 0���Wo����y��������V�::۰��S�qD�H_Ger?������:a;��Sߑ[�ylaNH�މ�^����7&��{�_M�.��U4p�$�V�9X.�ݷ�q�sf«.'�S�N�s�xJiG�X"Ͷ�"d8o��T7�$���8a���唵��_P,�I,0_�ߍR�Z}1�v=e�������	�j�:ؚ�A'ʷ�.:�˨-0�w�H��#��Jn	46�"/!�)�i#�Aﭭ=(d�ӖT+�i���Y~5;�_�-ldO���9��	��	A/9�|ձ�P9����f^G�.�:�,�a��<ަ�G�K�j�i�l��<������bXj����9A.T &ۅr2V�N�J�H,����bRr��tR�Ù*l>�r �b��"D�J�b6�Y�c['j�2D���U�8L�1����v9�:n��;�JP[S�q�9�+"�զ�D�L�����g��
�)Z���]7����˲IҔY�e���M��|��~q�6�_c�/,�����P�wW���)�aj�GD4�<��� �M��π��z0��Y��ө�%��wj%�"-��EI~��t��H<,?���!ȓ (9���h������\��"a���H�/�+��&���|�"�@'��-�7�Y���[B�a���В4h�Q���
�/��.�ό�Oڋ�PrQ
�ZM�-P?��M=s�2�=ô!��_)	�-s�dW�ĩI��3��H�A�mY����QQ<�P
k��sҔA��-��Ɉ�E)�'�5��.��M]`5F٢U�3nMz�Ww���Z)]?�Iy�V5MR2�
s��\���؇�\���l �d4RӚ�E"y2B90�mz��V4���xu9�������ۮ�#�Zb_����
�sFP�͸i6���%��z>���:�F���9�A)o� v*a8��hW���'z��C��zh���FNWY6h��a|~�b9��b.�Vͅ�J�7��
����lґ�Rh��e�\�h��S7(�W�"�!�
	!��u��;�˅b���7�����.�>�"�G7#v�u�&��V�<w =�f#6{х�?2���ꆸ�,���Q��"qL�������1�4�&=��=U'K��,O	�˃�$���d���K|�)�-�v�E�@�}ط*sB(~U�M5%��� E
NbQ�('ty�s�O�(��QݧRc�P�w��t�`���j]��R���+������ x�MR���?�ʨ=1�ħ��J%\�.������G9� ��V0�G��'=橴��jT�Ad��u��s�f�u�=_	-������Q��Ľ�7�r��
4�p�!�Ơ^��6!��.+$�`��3��r�k���!قIK:�g�����4|u��֗�R"�e��1_l���6�y����pg��ف3�������M9���Y��'�U��[��ڑNBȷ�2���i�~�x���	���gWS��p$�� ��Y5��s�p�1,<i�SKo��U�if[ǽ����Ƒ��Ȱ'VM��Ѡ�os�%��6񙎦���*�N~�9!��f/}����ݷ�"��?�
r��o��BO��}YS)��G5�����P����l]��%vn�284{>�E}xZ�^(���+T�
J�q�s���ڤ*��8��:\�XN���]��m/�iR���U(Y#�>L�=-"�X#aK)VChj�R�'=7/0ƈF�B7�w�j;��s�zi�(�#��5�H��ӂ�ل�r���Jʞ��Hx��D��,�p��0��}�K��DB�?�-/WG9��o���6Ҵ�>���_��/0�H����5��y�/��_��z��7�褸��..,�<�w-�	�����Q�,W��ڇ�͋���<����k_��\e���G�;�1�m�
Y�X ��q�j����04vi&�&F�Y,���]�,c`�7�	�?)���������	�0�T���nJ⽬��������b{L�� B���lU�%a��[�~ <K@�&����ylJ.���:��d�АH� ��W�D;�=)�	Ի)���}���YQ��pL���*���9�*٘c� �1�k:�%��^�o�%�&�7f?8Ne���Lu}鼌�&zH�!6�6�7̢�X��>�9�+�бxX�^�$��R�W	!��0+���Fh�ª�N��j.oF|��lwO�l���Ȯۮ>��U)�<f&�â�N�^�>un2�h�uG��`��]����tc����V�a�j���h ��"[\����
y�3�o䵌�	Y�mK�Lr���6[��p*幻N�����#\k�u�Qv��Ks��ςhQ�g�9�A�!��t0�u	`<�<�*�X�O�#J,���%��#���b�q%�� ��ᦩa��o�	�������9G��Mrn�'�" �ƵQ������]�p�.N�9�^v��6L})��������㫝g{8�w��H�wG�gD�>�ne����]�]��ݮO��nP�Ͻw��5�a�0���R�Oh��I�uN*a�!�*�����__P��!vsB1��£Z6�&�9;_��Ra�s�l���C�����ϣW3�z�n���ϋO�&�h9�=�7�tY��3hN��}�y`VO�f�l A�P�}�aDE���7�bq��4�k�F�WƆ�߼w�2�Wf���&T����/��/E
�:�떰�싊���ž%��F2S�s��C����@�>ƋMU���\������j�r�h��"ː�k�,^[�>�Š�h��������}�̓��Z�&���/��M�~x�kLf�t��2�>�)��n�?_�)��c��|��_�64u���Їro�\����a3�Tp��&��,J���m�Mf%bzZ���
��8]�o��Q����d�~,آ��j%�	.��^Q�tGԆ��������INX?>���s���7�����؎>���
#k �6^ߒǟ;ߍ�AI�b�	�[@}������^Bb���_����hIW;���J�1��T��P�ur5	�?v��->w��'��A�6�-�xB�	�b"�&}r\j��?3�@˥��j�aFqvA��a�Uڏ���6�Dv��P��p!�R��]&�z
*ڤc�t�=mƛ܁��"ؚ0�� ��:X�o���#�t�)�:��^a�V u`�&	#���<{�L�
?��=	��;����yD�=@�8k�Ӈ?���s���F{��)8B&8c{�������>��Hϥ凹�
 ��w��"{���a:� Lg/g7^���vk��4z����R�K�r��<�h�H���ޟG�R�%S3ӆ�b_�T3���[J�M�V%�?�>{�;ݡԿ7� �E;z�(�
�Z�-BR����Ԏ���:
�OQ$a������(��q�X�'�xRn׋��j2�h+~=�,+"�К�\���v�|�4���r�^�+�����B7J�}7ҒefJ t�_�J��$�&2LM�v�z��P�}�Q�)�ϗbm5�Ѽ��%���f��Y4N�	Z�ഐeTY�����HPʺ���+Ao �	��$h$��($���/��s��$��UHs�+P��Gi��¥����p*��)����Ѝ��r�	�cۑŁv�&l
�x���Ah �/t��A5(ճ�]'���~c������.+��1.�2IJ�h'��)����>�4������U6*�kX��D%WVbR"�F�5ۉ����l����j���L��ل�mR����h�o.Z-F2S%7�o=��X�(�4R�K�-��ȴQ$��	��=G8��zuI�S�9��o�f`E����Q�z.%��ԨP[��8� ��,X_*9�x��1�kF��yJ")��iԛ�6#f�����6��'��E�(�?@�W!��@������#)�m��.���,�i���bw��d����Ϫ�Ý�:M�-4��?���2��}v)���'VZW�
T�lۍ��A'^���q�0._�4�&i�^��|i:���w�w�^c;���{�Iv�y�vk\�j"l�G��m_M�T�O����Y���:餟�C��&�;?�!L�^1����!����'`?9t���Bl�,�F�����L��ҭ�Ȯ���X���ض�j0��'�S�m,�RIÍ�	v�+g&��@&W����f��(�>t	<�[�}\\�;9�j����{䁔 0V�S�7��.�B�9×M�Y8:�`�J���xr��f�|��Ǜhg�q����G���<�~�,�yrQ�6���`�#�U8,���f �9�����\�B�?�[��SѼ�U���1���$#V��񏟵{H�3P�y�Q�1��� x��Ӌ���"�������N3B�<�^�q~����ʣ/ �ꃑ�,^�O�	ψ�x��m ��Q�{8sRفA���1L�9|QP/p>6�K/��n0�2d�@ٱk�K��:�k���I�tӑ�^?̮p���ڼ�]=�_Ɓ����q���9}��f���a2��B�?� �ɫ�]l�� �8[r�	D��)o�K]�V��ϋ8���Y�[t�:�EZ�y��Th*J�ri8<bA���q���#1M�O������+0�l${5f�=v��L�
����f{a�[��.�:p)�O���S��S�|��[OC�Tw�ur�i���p�5[S�Vy��O����%C9
�c�(�4B�>G��S�L��p�V��>�� 1���)�ڜv����H��1�-��¨F�!P�Z�/��cL����D�f�o��OlL|g�~a�ګ�B�@2�ΙI�G3̌4&%�t��թ���D��>\z�,"�u��k:��Ԇye�v<�2��E"���W��P��� �d|����1���k�z8Se`R
׾;�2�
�O��ؿ�#iVm��ٺW���F��J����e�eVWaT]����e�®5�^)Ʋhx�f��"	��l�=IY�o��j�dY������_#�s�$��>��js�Ah���3�C�k�>�y�H����$���m![e-��S}t��M���W�����L�VE����! ?3$	"�������k}8�}ے�9�Kx��-��a.��ބ�jԐF��������Ql�;!��7ե/:���>*s.L�M�H&ȭM����t�-f�k�0�4h��h��i�q	d`R*����~%�ߴn�%$o�c���"i8<|��.$�LE���������dB<��i;�/���P#>B��pbb|�9���6%��\:;a��e�#k�hySP����#�}�o�溞�j0�r2����"Qm|��&�u��,��fŖ���S<�~?��W��e�r��t��bF�����	]�ϵ�z���N_��e�r~�o��$xٜ݈A��]wc����|��}��{�8E�tT�<�Zme�)3��$2��t$����->+�9	��uwK�g+3�E(���q(w	_L�����H8G�j�`��C�n�`t�Ў�uay�PXh��LY���d����v����(#��w��X�^�� �o��T�I�\�}�@�	������>���ؕQ.�bk6�$Mu��q<����b?<7� i�W���W˝j��|���T�A{���T�e���N�~%�m}�4n��tw��+���:t��I��aJ�r�~60�^kƲ�o6�ff�]����6���aЅɆ���������m����m;�"Q/ ;tg�%ӯ� ��_�~I���2�Wsy[#�D\x�����hhFzUwj����e������hL�Y���#kY�3������N�t���@��052@pl"8VE������kW���'7����m��;FE?� ~�����-Ip��>2
;�26t�9
PxQ��5��L�,�Wh�*��������I�rs&v<�*>dq����	��Zg`ܐ��>v���c3����E<�ӆ)~�4�(k�-�I��϶��r1�<y.�����hB���)2f����6�e~�=�V��*��pb�d�fԠ:�5v`1�nX��n'>)ŧ&�"ZZ��t�J�D�����,k�����T��~�7$"�8��;G1���'K��&�\:1�d��E@����G��ڨ@
ȾL���p&��V���q�"4�\O��lC�\N��85IAbɞp���)2oq��`��e26ކ-Փ��x����Lo�^� O�WKqz"b��Z撚W��y�4�p9�jr��>D��2�}�w�<�qou2<���<l�o}(^��.�9�M+����&�ų�"�|��_c�`��P4�Z��f�V�4��B5���7Y���$)��w��_%�O�`ཟ�iz|G� ���[�e�Y>ّ�Y�\�^�0v30�p�>B u?���Y��͗�s�����sD���6�3q�n�{;��X~)��;��b���1�M �<6�G�j@�iu�S�w>��15i�i�����j-�~���R�����+�s��2M��a�����S^�N���L�����`V%F|a�`�g�E� �n�Wq"�׌"/�� L�Hd3@s���αA	<@L��E�o�sp�} k��x I?r��o<����F��9%0n3���	Qn���;��ɋYtzi����}K�!�Ť��M��n [���hx $�E�	�!����}B����M�q�7,�p�hZ��*���KU�<V�Ջɓ5)�m��F�E*[Ә�.Z��q2_]j���߳��$�[��+�PH#�نz-Ik��
X�I��7���JXz~���'��Y�%�<r�F��'�"Tr�J#�[��<�����T�Ը�F"���_���eڽN!4����5P��@���.���	��G��H6��h�0�!ȉ;#��J�u0'JQ�ۀ�l�w� �<,�.Q�
䀾䐜l!��M�}ʃI�?�L��׷�\�N��㐿?T���*� * ���e�Z��҇�́��"hv�!�+p5��P[�[��qp� P������9��6��k��Vc�TX�y��6:̲�amR������3
��=��o�췹�"����w�$�RS�d�K+w�����&��5U3Y��ha)�w��m�}�T����Z
N���/�43�3����+{
�nҘ��"m6e�9H�F��-��\�d���U�D�57��P��xkf�����9�4���`?�M�IIT���컭H����憻EEE���3��z�r�W8|�8�\�9֘����� 	�s�W@�@�HN�-��t�¯̌H�,����@���@�(؃��p�?^U��5(a,C�6�~��vδ:5���E`���.�Aj��Y��"�����!x�7*�UD��
�ˬ[7�
^�D�}��y���j�u �'������Dw�ݲ�!�!�<���ͯF���.X��]�v�(��A�,�g�=���e�uN��I���$%�/3/T�?�:X(~a����m�ܣ|C���vK��W�R/��?��2�$�[�3U��xs�j���k.� ػ0���Mt2qT�N�m�[�.V�ݬ[��ò�}�����ݰKO�tn\U���9Y�����Y˸�#n~f�G�\��1����3s��I-�e�2l�,��ԯw�ʭj�5�m�g^�/�����"�b��`�E�ۅdT��uA�r��U��u�W#Cs;B%�{j��建�Np�� �Ӿ�?����i���I.�qPCT�*ȿY�J�H�Py��c�% 0ހa���0���K�6M̠6� x/�̋���V/��S&�2�&���bڈ�q
��.�j�$L�J�b�p������X7�_Ư2`��_��6��.9u��&��}���he��6e��>#1/D��9bn��[��ʪ�q=��Kx�ǡH�۫j�����#���{GL��V~���{���
�T�!���\�޲��ֈ�̔�az�6���ϩU��ǯ��5���H�Ͱ�	��n�b{�+������E*�^��n�Lg���y7�t7}������,|���zm*� 7v���P h)l�"0�-������n��	�� _X�y������m��Hkuj:D��\��N[R<����������n'fh��k�֥�wW�D�V�st��E�"���gm�L�/�#B̓��,�i) ��._��EhL>�����:��wޤL�R��忂�߁��F[G�XB}9�)��/��,`�m���dl��",L6xhL�ޕå�
�>�++0��9 ���7���6i>�L�����τE9Y�b_�X/���~�<�I�|y�n�n��q5RR+d��ǲ9�79�ԗ�:C��J�)��<d��2�3K)�	1�ɋ9�|(gg��tjA}���臝U�nq�����#4�J/4'�
-�9a�AI����dũ�%����=�F��q�r@,��x7r�v�zhX3��fڒ���*�y��\��N_"�+�� ��#��C����r�+������s2�yS�iŭ3����U�<�d�v(�\}E����~��������/�]���K �|��X��'R�O2�u�����XO�R���oܤ��=�W��]>:�N�j~�:����2% �j�a��2��q���	Ҝ4�!�{��A[���]�Q_+��>�O�����%`��*dߎ
�X��l�nN�*C3~I}�� _�)hᴡ�ृ�,�R�Cq}�C�������w�,6��kx-�ϲ��OJkM%�9��.�������MT��n����i3K;\����SV��@��܃q���klk��+~"J�����+��Ӥ	���;�=+���q
pvm���L��%ep_gv�W3t�G�}������`��ES�5P��̾�YN�7r���n٬��6�uqXS�u�a��8:ր4������Z�k�]���Vǖ���&�<�F���x�ؕ~�$�Ӈ ~x��UY|��}<5�����˜��u���Y�lG�[R�ܸtPr-���M'ך:�!��^r�;��m[X��;͐5�v;�S�ܪ�e�>$yF��JK\p���k����R�e`��ˀ�:_3.���\3rʭ������"��bx�)��س��˘��%*tT��}���4mS�'�#���r�_��<�5.�ޕW×Ɣ���D����(#��;i|��8|Q���ٶ�|,EAF��H6��e�a���F�A�!of� }Ap N��58ʶݤN�e&`���?F���U�)����SQ�2�,����S� �$-�8Ұ���w�t`:�{��p�f�e���a�`hgG�k���,�s���E�E46.ZqV8�Zϫ">�D}�
��2(�S/l��{��W� ���C��m9W��e�e��u+$5`�Ó|�Pu=�n��n��Y�/���rD5�I���h$aEX���?���3��.y͂!~֒��r!@Bz=�M��^�Zl���`��D�F:o" ����n�x����#y2:�.������Bf"ҥ���R>��ckA�vֱ<��{ט���N�t�Кf�S��U�x}S���f�nٟ�b8;�J��|�(�v�y	Ȣ<�;z�X�U��������i�V��^a�xט�����E�  Kz����s�b�-	 6�����U����dQ��wFO�l1��](�r�R9��t~��F��	�0�}or�x��u�Xyҡ\I[��"�AT�0cbж��w0_�A�H�V
-#ϛr�����Ǖ�:�"(S^�e��b5������X\Tw���f��mLxT�`2�#�,�[`] M3%.1ǃ��>�K�&
�d��E�'��8Id�&�.�譲�Q���g�@��Yx�s���.�J��4�*�D�/^�S�q\���3[���NU����R���8�-�@��K�^�_�F�ڹ��!��a�G׾nB����77T�N�ҁ�q"�@d#����R��y����Y����d�b�j;79P�f��??�4�sV]��;���%�d�V�S�cO��U�\�������	�w0�5�D"Y���aM<JӛI/ �����]"�ˆ�,��U���]E�0e8���q���2�5��I{b�Y���K�q&���U��+Nk$j��ft��gG�r^����Ņ�wЗEƋd�����:I*7J�94�m����ONoB�V,=�&Jf'JeJr�~��g�6䝬�9j��r�;��J��0���k�'���{��p��Mė)�<tLV�q��,��gu�<��;ٛ�C0��"hَ����	,^C���ct�,C{p8��Hv�gE7�Ԏ��A \2�	�T�a�F����ql�],����� ��ۑ8E�>���!���e�{��Ub� Kc���xK�G,7"�%�=��?3���s�p�k��U5�<� (�Nf�3EѿM��|�C柃�z�qhe����$� E]	�oE��Q��>g��B'ae�8-R����J��#�8@?I�\X�9n�7��0����k,N�#����L�lpvl�������'�=o�QZj�{�%9�����9P)��$�f)A�)}6|�4i����%:�R��'�i���͡��'x_�&��N�2_o�{V��y��������7sZ��p�$�x�$H��\������Y�XQ���^/�n�!v6��dL��t7�}!d�%.��Vf��pP�bĆ:'Ҫe��u���P'}�'��7G�s]�A�D4>;��D@�w %���Bt&���d4�T��j#9.`�,��B�EZ�>gr�+l�:ا�������r:��َ��&�q�Q��@�a����s���gYiV�>Fi��ؐ�P���h�WA�����= fc�����Cm9'�+�x͆�SH�
�0Đ���yr5H�1�~��:"&�y~]�7�P"�H�Q�?�BO���B ��e:ؚ�Uo�qs3��գNsU�Gi��{I{�6���9
�m3P9k�a�������.��h��Ђ�����i����������^�e�YS��.�-}�pt������;�g�k���6D^�5U"��D 
�˚�� �B,�6�@���m��&z�ǿ/S�+��r&����I�ы],���S��H�T���n`�S�u���O:�dV���;#KTx��z_,�5�0��ɨf%l�w�l�P���gi��O��D7��	"��yS^=�r����E���Y����t��RՅ�4�&_ka@���kls��V>�SZ�wX�(����KZ�W�_��^$�S;R�Qb��:��ʙ~�^ �Y��7��':<+^Zt�~�����v��㢧߶Xa�~���z�<2������^bG���w$*S,:Q��Ľ�i�D�dZ~ˁ͙ϴ��9�R�vi�r�l�e)�c��J$��@=K�2%ݪp���ڦ���y'�l�ْ�Jd089����Sc%o��,�@�ߘ���}���C������8�>�{i�M:�o�5䫝������T�0����� U!�v���[�Y�����"�pҒW 9�{���pG��������Q�6/a�!�mʾ��3㓤�-��5R0|$�
+�q���Y�-?1d%������O���<��pT�o��M�-�IwUs\ղ��,�F���l��5{r�~\Q��	4S���L�#��\.h�%�.Y�TK���Q$N^I7��?e��]1B}�]
	>�ߟ>�=���>����c�"�G�yh<"�G�l��ܬ}��p
p��R�����C}]L���6c#?��j�R�v�U?,9 n�1)���|d{#��W���W���=�4I����*���:�/j���
�G�?� �SA��r
�;\��.Dw�ބ��-�$�َ�ܣ!Z��/�|U��v;7^c͌,��0�%��q�.��a��ު%���_1�SH�	E��e}Ŋ�=w?h�G�߅q�_���үE��udP[SUY6��}y�����>B��d��A\�����f�x���qU1sz���xǔ��q�Z�������P�ϵ��F���a� �RJ{��֚B��%�S(�e�_�i���"[U�orW�w�K�U���@/�Ƣ<�ŭ�t�a�BQ���E�A��k.�������ow�s�F�BO#��ԥ����e$��?+0�~�dyծ�}].(Κˤ���w�7T"'`��V�/f�T *��A�l�{�0���ߝ�!�v7h�sAPh���c�,�tKzIZ�c���f��YG��ݴ8KZ�5&:�i{q7�X��'9�L�`!x��"����N��=y���_����z�P'�Z�������0�3����X�����l*�ZPW�3�d�ʕkO�bm6�Z'����^�Y�5r>��ޞML����`��U�~?�ّK��	�r;�%�<�C%�J+ȚBun�:kl�fB�t���2q� =�K�
�BQy�sѶ�&4*�vw���6�#E��	���{�?o5�H�ci��٩���P��N��((�fN�F����T"��,H��v��cN��p�k�
��0����_��tXfiF
OvZ�q��O|_"�'�Ve�����fz�S�%�14`+���j0p��F�?�+��������+�rw�pVMg�^�XR�/v�1�[�h*s�?<���u�y	p[K�и�Қ)zc�8U�|v�_Y�*��֭�ɩ�ZU   ����7.<r.����G�fۭe�"��}�������؋���OI\�� ��G��������w�R� ���7�� n.�YS�,J��,@�>�þ��!aV��F���-�k��K��_ǡd_}����Ԇ��$����9�C8	�+�Y�V��30T�>L�`-���v���(\�0�n[&)��w��z|F����ղVUIze������࢘��
:���͝��<⯢�3�;�=����;���AWv�ꞟϦYi6Y���������7���K��zEU��)+%�]�����dd+1���Ít����H
#G��d�i��(H���%�휁g�4Lz�U���^�!�c�?Z�yis�lx�Z���-��M�P���	t��j�)�� f��2��_:�v<d��%S�~�m�FX'��+
���]O��W��/=<���u*�خ��Q(o`���;�wz����<��f���K6�\�(� �O��+Rzh�C_f�����|��gf:4��'���*;7��ś�G[��q�,홸k�su���܁�[�6�B5<�zCЬH҉yr"Gn���S�:� '�8w��$~q�sn ��z���X���PD����At�r�� ����9tYN]�7��ӵ���(}Z��+
R"UqYC���H��pF��,kd�NS�t���z"���/PҪ�jZ7V�Rh�(�H�4̬��UW���c��]O;�ؾ�pV˭���=��o��Ƨ!�4���q��*ƛ:�tfמ(���5������ˇ�\I��ʆ�F��Dc��_4��Ζ��$̜%u+h���A�c��O�o��(:#M�$�����^yѯLa�5�K����\�l�='�Lh%b���,��9�G��gz��v�|��h�a�:�^	W�*,��s���ݺ� �-}H��	'�%r`+��ں���4Ͽ�I'�-t���]�_4���Q�ZUOW� �^F��Z��B�3��L(}����h�a�]!�/Њ��n/d�G���]��lϠ�x̧a()��:L?�bu\;��h#�33H���@²�P�Mb���E��'�r����|�!k�=��y��/�xr"�?؆��?� ��זW%�����?�cu\�����Xg��� �,z' Ԧ58��|G�m�K�����t'u~����8�sP�7Y%�nAvЂ�L�1�c�_?2}�u>������8Ra%���~�	]�Kcp*�1P�`х%>�Ă���r��p.�K��|�R��������:���3��zoUaN��LQ�����J�%ϒ�*�@�SZ@~�t�H6#��&8'��+���/VSL
E(w�egpk�
������t��.ƣ-@��UB��P�8(��G��|:\)]GjJ#�;dOjm��]��/e"��gD<Gʳ��0����<y:��;	���E��M�v��=Pi���2�l�`�	��U��ԃęs�ER��DB{kB׫�*�U �4Ye-R���Yk�!��҇�_P��Z��Oeó�ӺR��Ǧ#Z~�E�]/�7����R��H$��;�Lx���Q��N�4u�b6m��ʺ�~>�6�#���'�M^&��Q���O�"�|�ȶ;���1S4��r��ye,c
�X��	��ߢ~�{����:N�`�ц�1}o~�BJ#�$Rl����$;R-��OTK�|���A���͌�'��������4f�&p�$W�L�T�Ǧ������n�и3�g5���;�[F��12�H9?/w�`����3>{^��f��&�O8
Zo"	�%&��_/R(~�_��e����{'s�5b|ߤ|fu���z��W:{�/�*P�"Dľ8�>A�%Ri��u�"TԟW%Q���u���VP*cd���)��q0x�!�=�`@I�>H�(6�N�����Ňz��pE�X<K1������F�R����!�{������ [i�x���4��C�v��>I�{�qn!��6�1��
Ɋ�
�������B_�y�!!�*��e�,=�l���co���i5:'�L�]�b{�t_�](o��ד\#����o[�[K?�H��V���	΄��~��WSR��9/!_ೞ�Ԍ<��/��>ڗ�!�Q��o��]"4Y�_ި��!�������̄?G
�=���oh��¡�㷾4�P5M�8��B�����'��gw�7�U���!&�\_��Ԉv|h?M��)Z+> ���e�U `���聹�V%n�]�$m;&�e�=�\�����SD^0a�2FLq͖�v�z��Z��m,q�7��>�/X
�!/�QW �?*ù�$	�+�秕�Y���`��Q�Z�E#��/�O��X��X�����s�J��-Tk�gl24ǔ����UC�U@�?0Vа.��s�1bԜn������4�E������O.��,Q����gW1�@��f��F�����Q"�ب����/ʵ��a;���T~�9�G��9�,�WD��Ⱥڥ�W@�o�qUH@j�(��x᳞�=Z�R1������MU/�Z�叾ʹ��FP�h�(�[��o�'lF���Չ�6�3��� �Q�,>Q�Pc�]
�j��U���6ܤ�1Ҭ�C�y3!K:M�@�!���#Q��,C�� G՜��Q�F��l���c
c)f���h����g�-y_���G��N;��F��|~�1fM1)�����_]L���� M�+艩[ �K?	䣎�o�rf$�GD���������{ؤx��P����1���!��|_']껡��.�����Z��՝�H��� Cg}�>�y�#��sQ��>��S��D�D$�P�@)��e�C��w��y�'|JE2J�k-��G�����r�s����h�?0���lA����o�Ë�U�yn�&�댟��?��?��p�t�s�+IƎ�o�y:�����&r��S���ixo��U)�$��]��l�Y�3qk$�_x,�aOr+�jPu���=5	G�4���P
R�;� d��V÷�S�(��&f�_">G��O�@�q���²a63���A��4K�����k<	F�
E*��UԢ�ҟ��(�;��_:^��h`��^�y5ך�c�=��\)���9����S6v�ƌD����Ͽ���D���8���(��b��&�62k�Ҥ���X|��h-p 1�Z�����J5�fG5���N�_{ݜ�*�����@WM����T�ݭw����nW��6�}���;r9`܍�ߎ��Z�)c�ʆ��à}�=m`��t�����6[u{Pb:p�:ܕw��FF E˱m+M�=��=��J��_�{�0��H�	h����m`�]��08v������ޥIK)XM�i~l%�4U��$���2�dI�pOV~��&c���ph(��_��x�L���g�Y	�M�$5v��0n�'8��
��#@A5�J�1Ȼ��n�[�=*-w�kۙ�`Z4����E�I��m]�9R~��WZ s�<�^3����/��`�u �t��B�G�v�����������L��g��Tڀ�͈�o��$�z�Aţ���1��?L���u�R��g;w�dm�:g�
�ߚŀ�A�7"��YpZ��j�?�����`��������p��]q���Wn+�῅Ĳ�L��ph�Z.M8t6k��$�6�Z�[�E�XS �����c�n!&	�ְ������;5����EP>�;p�h�DW��|!���;�Gs�ga$�;�Ig�̫�����_]9,<�g�u�T9��lm(M�A!zph����՘���_U���@�����MNiW������ܝ&	Y�I�����W��lZ��F�V/��$�zCl��P��~ �1f�t$���Kh��,�b�z��z��Tl�`��'�.��.�&`�D$<�Ol�u*�2jE-́�#0���j��&�&�|3�i�K�榆���c�.�64΂"��!5ņ�M�����"�j���uM�P���s㻬�|�TE+:���6-J^1��V�B��y蚼yԘlv��z��Z�d���cH�K������7K�����?;�9*�%�n�"���_��
?W�d���/m6�y��=�5�?�asY�3���&wNN���B���U��nv�}�eV�c����P'9نsj��M����`�s~��f��w�ӆ��RҼ�^��c�ܙ�B����J*��zjr~�C���#Y�aJ1��-AC��;I6��t���-�j%�g��,h9�'���Q�
�G�7�h]��5�p�=�P��%�-\�V�[C�½*�$KLf`L���lł��a�W��O!�]�HaY )#*�t�֖�>�l��u՝����Zt!�q��á/-��[�J�sJA�>ϙ3&7(Q��d��T#:I ���\��ր�x����Q��F%�Ym���i���ax,�S�5���0��3�Ks���X�6&�T/�xb]kw��d�.=�[���<������K��$��>�V�ī<+#@˧5����_���@��Sd3v`�;��/\W�s;�)�s�"w���jy����g��p�ՖH��w!>�\YP�(�tM���`�$�/b>Dv�߭�ݰ�W`u���RvɆ?#�N�%ؑ���X��hsL�T5:eG�*!��ݺo�K#>����ۨ��"�bW���m��[Su�m�b�S1)�}G2��s/��,�gx�����5�,�����Uf+��꽇��C���g��P/&%���N�u2�¢�,�\���qYV`w�د�Xu �u����-)���˂�sy+�m-��4�E��D,�	!���NTѦ8�