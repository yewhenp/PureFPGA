��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_�}ܛ��.��i�F~�~{�J��C�a��K-?�<�>y���yewY�&�_��wr��� jK���w��C�Hxj� ۞�
P�D
��6⼞-E!F8��ؤ�Ct"�<&���H�����v8��#��B����,w���S�T�Aw��8�ZJ�*K���,3�3W�݄!�Ā���ԕ������[]7Tguб&!���t��R7��k�t��@��atUOx��1ѓ_���T�g���c��Cj5�X��53��\�S�(�E������fS#7���|�b}��P��P�^lS,"m5j�B���/�'�0�r·zv���}��'^��.5<{�ەw!4�/כ��޲�a�ŝ��ݡ_�R�LވG�ڄ?��<��3��
�������LM�T�8Eb��Gz�"A���������ռ	�s-G[)B� 
�\rb�Fr��{��q���J5�^�g�4��ϳ�I�� =p=s������OM�:�K��]&�j�8�v��W��k�������E���)c��!>� ed+v ��IW1�;�ĮA����.L1�Ξ���"b}�9�xe�3l��������Ƶ��ߓdf�m_����ҽJH��|x/4��q�eMh	!T���|���?]�_KU���g����{x?�B�T�+�%��)l03X�I��iHE,��2s��<AM=����5f�pJ@q�V�s}����74Ws;�
��Ti,�KJ����p!�B�DI?~�h��N2�T+EMQvq�&v3��TT�ͅ�-Dw�����e7hZ庳��5�9��=�b���02��$,������Ғ{#�^�w���ִ��=�V���%!�	�.��/<�7�0��|�S�1n7&Ι�]m8�`�.)��ֺ�ws�(N�h��\�|{I��M���&���%��I��mO�M�.��<�Y��CE����3p�n���ҭ��ɓ��U��<�t�?6
m6r�i8���g�F/^6��ą�=E�B8H]�ŔӠ:uv�궆3P����X�XD+����qn���u�3��� ��<^��}�i�-~ϊ�LG�|&沀�b�Y95h|�{��u�;�H�	l�)�dV�1蕫JQ��l�A� ������$!����0`b��6��j�@I���M%M���}؅#pƀ�}�Y[�o���ݶ����|���A�^�Ž��r7�+/�������Y_����p������I����3���(��	s4�����c:�4�`�T�SdI���)/��tz)���Ϗے�N�x�q�����:�ѱ�Bw�c|�m�	۱
[�3t�!��'�Y��U<U�\i�NV|���u|-P #W���Y�1�R�D�uc��FQ���d >�g%�����s��2��Q,�a���&�ۃ|���L����R��`U�a�O�G��l����ID^����iݯ[,o=�
ܷB
a5OB�}��z�?���g���Tz��Ͷ��A/� �v�T�F�����E�n���H1:�g��V��'�
�r_��s��Ho�ݘP6`�����ЭE�$"�RV��ѭb�*ׂ�X'7�^( ��kH�P�z������S(��H��q�1R��¤�DF�+��Ys�ᚏ�$�N��)gV#�K<@㉴ƕ�.�c`��R�>F�����z1Z9h�����=�UDG+�/c tv 7>��f-q�t�ο.�4=�� �+}�7��[��e��mzy��P�1��C	P���bS�K�f(�z6��q�z����P<����\�D���d�o�q�fN<�	/Z��T&��EP��A�;Y��zu��MD[4�HN�[z�q	���u�������,0�g�GX���:���$s>�?n�Z�����k<�qfx�e���(j����l��<��{,��m�4dħ�Sj��/�'��;'>����S����a����<� ��ƚZ�5��-��%���_yh�y�� 9���y�����?*������	A�� ?�n�0�`�Z&m��.#B���׊�͹k��Rph�|��p����Ջ��rHx?���T�*e�
J4�f�	]3�M��cAf���,�P��>�d,K�BDR�J��+Jy���$X�s.���'�^�|����*����&$?�ڸ�E����[�N���:̪�LSU�M��m���pW�����#h��� T� �����~�&��e��wN���m�J�, T�9[.cg��2Ä�g�����T�PxIw�[Z�Λo�I^ޓY	g�&j�
�,�
�������Ѫ�W}���Tr�(lv�v�ɪ����XF�3I q .j�O��[]�t> ����r�$��閛?� ����65�|X^q��c��3��C|�/v��'���������Iwc�|��v��{�䠣�r8}!��|�����:`0	�����*��:)��:跕p�$[�ft�Fc�v�q9�Z����S�v��ݺ�s>3�oԍ�y��x�'f>^Pj�7 ��rP�Εx �S��>���*Ԗd
��b+X�]����8��??Zj���h��^���a��K@`O�}�nc/қ��J�i�i6��d�!ķ�/����!�;m�V�U�͟��"Lj��24���k�Xm��w�@�N�tq��~F�p�[���핼���ӏ;a�d�p��d䯫wj��Cb�nM>G=��pDB�b�=�+����=t��>����A�t�tq��_� N!f�F$9n�w%�W2Ә�FHXj��YzR
�Z�֍^��=�����n�1vb~�&@�̹�é}���h�)voy�%�������L�^�����pa'�2���"ϵj��1L�1v4����ڧ���t����A<M��m0�g�ʵ��@O��_��=�= ~�b�U5�N�?t�ye�F��#j�� ?�lb��u���T㿄��۰��t�w��{���a�I�WPL��#�$g�]v���2x��!j�/W��0��JY��m�g=G��m�5�Z�0G��A�OnÄ́V�$�Z0�u�����	����\��5���U����6���ǁ*#�/d��[�s>�~}�#�6�L�@��kKAɶjeB&���nVO���bz�l��L
z	��������F��1t"���ӹ��l#��Pz�϶�ɫ��'�2(w�cR?jaf��%���Ӿ����g��f>(a��z��y��7�@X΄�?u� ���;�خ�Dvwhz��P�	8E|"H��r�7��*[�X��on*H� 2#3z1X�fP��A������z����n�Ԃ��`��#�r�Ap��i�=ťi+�ː!�y;;lTqk�=K$]���%-�/&�wT�~
q/�IE_9����ĔfA���ѵ��������������rx�/�ѓ:/�C`�l�6�*�sD��L��=EUä'�'n��	UQK�AR�'�u*�]�A &Q*��_������v^P)?^a+����>�"B�?���¦�����n�����֢y��,�A��`����Z��sv�%��*��ɉ�8����'�"�T�p18��-�o=%�Yx�WK�X�_L�������M'F�+����dK��N_*|)ֹU�`���Sî��Q�/Z�}�;%0�F����f@�C;���g���iQ,�$(&�#�Ŵ!�NHM�P
ڞׇrO�6e��	<k����g3P^�[^��i��Vr4v�~3�*�	��39�̮� y���/��c�
�c����Շ�(W�YQ\d��x7 ��i������/l%$mƷUs���FΗ��a苦6�!F��\�ʳ�ri�hZ�H�6����mz|�lz�g��8���`��j�ʝ�O)�k�����D��|{`s<�P�N@j��c���>s�4��R��D
ĕG�ߊ�-��db�*F0�=]U�Ml ��u<��c��|�!nPc�O�]�D�b:u��J�_�zj�V����)t���X���>��w�9�jk�
�UO�HE������H6�m����{�-��<P��s����$�-z�2FU�(�Nﵱ>�^=1K+/%�R�]��߇x�L ��߽H��a��Z���W���4e�7L�����R���c$b}�Q[n�P�>R�hU
��Y� �-�3B�e��N���d�� �nJ�Ѡ}'��=�Ɣ���$�SߩR32���31��9��*�Ŕ�t�gդGf!�@���NIqú�;�'m�ɭ���Z��W)�I�e�;�;���W��[[���[�^�
���s���S��L�:�L���ige��k��X���l.��ו�ȁ_QG�.����ټ�}#�px���8+ )�<�����3��JcN�X�Åxwb���j��o�ѩ�L���ʈ_q��  qD���:�/B�'(F�of���"�#�v�����lZE�K�&k���f����_�z,-&��}�Y�OQ��GX_Ǿƶ�+r���+ �&y��HY�Uy"�X�LD��ғ`�r��o*�e�?�v�kWr"]y�t��H�h�YzP�/��lݝ,��ͪ-�m��Z�5�<X����0�)N��#���ҏ�Hq���,B���'�avh�Z�b���~�;d
d�����������Z�r�.�Kz���k �c�� ����l�&��;4�����I9�� �_�a3{\��K��}���&}�$�Ѐ� Pp������4��/����}��!~�EϿ5�K���%�B��G�*$J6>֖��0���13�O�q]�B�xl|1N?���v��θ!mF$;`?��l�`4����a�\5&&J�1�1 ���59 �Q��������
�n���y�h��P���o� ����d��_��g����?��n5�U	��5B)�{+ـz5u}⻱*K7!c��Q�{Jt����f�z$�	���M������j@�-1a�]�]M�f�����u�����"�:f�s���%Q2�tS`(�74�Yx�?���������4����Ë��NR�鳏���n��ߪ�2r ����Q��^�����X���h�u"�ⅿ���T3��D'3���(py�\^F�K�J�t����Z$:����[���H6�͟5<�k%K�t��Uz�:��&e���-��<)�0^�")��q�+ i����h�kE�����Y+�	ό�}"B�3H�XHm�h�@�e��ܺ��*yñ�q����Cڲm��_|�0����O��_�9D�Ku���m�A�0-����6X��� 仪��q���-��t�$^�^��.t�֝W����w��T�~�BY���>[�ƷanM���-}�bt2���F��5$x��xР�`t�gP��I�AP�i�e&Z���(Vz�rTSb���QQ��Pc ����{R\+h���Qݟ�!_�1����1�\�}Ϳdāu�0ij�t2Kcn��	-ɕ�p:�p��uۜ��u�(�#!�3�Wz"�9��ǹ1`�N#j�)G��X��[���Z�j�\�Ś"��y������Aį�u=G��&�$��_��w��@�4x"�4��S+�L9P`�րl��9h`+їƨ �y�1.�ē� �(�a���N��y˗�<X8�?r��%����5ү�����΋l���n��n���2n���2������`�r1p*���Aa�`[{S�v��D[}Kq�G�"J|,�s~?ȵgJq�xB���0��F{޷h}��A/$���ŗѦ��`���J��x�����#:��AQ�Oı�U8L+�c�s����͡�g��P����{
����ɽmʔr��3"��n�pmq���͐�A����̼:��+Ղ��_EmY�0}��C�u��%a�+=W̅ؐ��7O+��2���Ը����{�͡{�<6@O*�|J�&�v�_ٗPU*+ �b>aR�9$.2[N"���k �E��B���׼���#i�dGx��>��2�rV�v���L�*ˡ�A�t�����?���"?>��$�h��E�C���kF��J�{����b��-�kY��=�)�mK0]s5��i*����s�� �ߣ�.U*�Gb�TS6#���t��*��!}=��h$�5�)���z�)�*�h�����ܱm� OzA/�9D��l�*��2�9c^l޺�c�c���̌��a������T9�Y�||��e*�	ʀ�/��]U�څ���(��Z���$c�^�yQ���a0����$�Ґ���tq�ܣ^����~WE�Ġ�t�m;��#��*5>gVwג�૨$�d���
\	g^�=�+e@�����]\,�e�<D\�`\
��v�s��a>���E)��\Tx���Y�(�C���Pr��uiY`.�r��5r�����^��Ky����o��M��L
7Q�t0 }�|-�����O������|�*�E+�������z�KF-Ԡ�N��%�O;e���$����xY����_�k�ۄx��T�~��
���d�7���=֩��1�//���Sh)��h�	��Φ~�g�8�cm��e�X��&���k��$�?xm�ӝ-���0�6aȇ��p���#�<����0�$�n(&��?2��`!&�gU�qA���-?\Ɯ�I̧b������v�Đ�"	�������v#�V�L��J��V姝��E�}�>07B�G��˩�|fb�K�sρ1l
�jsD4�v���66lLe.�����-�]#�I4�\��?����Q��E����d'��q�<e�EX���$�)ʅ?����r�8y�r�R��jiy^�H|h W'���N�r������u��V�ܚ������*�9���P�������\J"q֙% �o܂�׎�M��o�>���+k���ؘr+MZ�^6��B ���*�u�ӵx�o�6Fa[�N:m_�� J&�(_���&�669�o�<-ېU�
����lן������|'��_�ߟ��.���RM�5���9?���2L�[�`p'�W3_������YL�A��a���O�����/*��J�D6[M#!��0��^/����k��V�5w��.���F�-�?����HUC����ט��=.�C!�v;��c��)H.�`ʯ=km��⃅��A+z�3��в�h�X��.E5p�0dbX,�!G�+�h�t'�W��pt"q�3��<qm/��op�݊�d\#�����H����
B$����Gq!,�Z�I���l���V2rL�-���"�$�h/����'�����Rj�����$�OQ��㈚����TA��z:t���6*�p�՟ܿ� "�[�N���)��۵ը�M���vOu/}c������m�U�Z���������.'ҥ����k�3 �w�I�#anQy��_�F�p�k��t�p6�q��	)LŴ�p�����?��2���h�����v�����p'1�[�U<�:�{1���}8�sE93�˿֖�/v�� ��W���.3AI4��r�Kt�F���zH'�`e{�i�m�a�c�}
�O>~���V9�$��	(�*s�3�zt�~��17�(̑�|��ԟ��U��a~>~�B)�W�:�_ �k>J���J[�V�,d�Q$]�"��׈�)�(�H$<������4Y�����	*�G�8�;��ް1jO��|Jĸy�{At/�zsϞ "�x�kW�[�5ĒU�绮=jU�ָA�sw��B�mfecU�|�ܺ-�[^���blfn�.J|C���q������c�ĠN�A�O�$f�b��$\��S(v�ϣ���۟�3M~�I��
;xJ9�f�9r���"��,`η�U��������|�Z;/�/g���t�����we|�5 ��Z����K:U�
��BQj���Hw�o1 ,�&��8,Gg���ϻ^�A�i	{o�<Ӌk��3:�Rʞƀ5�x�����5�(����I�t�Yn
y���>��p0��}s�t��yp��K'n�xOz���%�h2������L���hKr)j/�G�M	� ��|XrΣf._�U��N��L5]��y�X�t���@v	��t��j��� ee�Iv+�^�j�82��,N�n�]'5��� � d�O"֔�S�0�_)�Z��!~N����kD�)�������������`y7Gd=br\(��p������'�a�$�"�cp*�y�Vn0$�V%��b>c�v��nl=S�q�5�A�w�Z�.�ڄ��B���8��8v�"�V�-�3@{Q��`��6��ѿ,��ìl��]^�:g��!��6���)5�z������]�O����f��(�A��B�~n��,UQo��#w�*�7�f���`�A2(z��H�`a�xS�[B���)5�6@�0��L+�W���V\ֳs`�`#�����+��b��9�P^��U׉��دt{�x�J~24ث� �T��]�!�Ѩr��k*�_�NL�lJ�^�ۭ@[�LF���)��=���.����>t!��A9�����ʏU��ո�(�V2�Lt���q�M�5���%"G)P��H���'Ǹ��y�y�p�n�n��dv��va�"�}���ǁ`GFl8i�|ҕ�r[,v�Ǥ�Il������:4�-̇��'�����x-M�P�+r�Y��ir��I<����j#��J�6_�7Y��9OɆ��d`�Ŵ��"o��w򬨤Sx������(�$P�b�!�#�ΰp���H!&o�ӷ��o�E>mb�X�)���M��K���n�F�W�D�/�П���i��1,s�Pjb?��m�(r-��R���Au��	Ք���jnw��%mlH�]�"�B��N�6�����Kh*2�Jx��\����.�˱��u2���)}�=P�	'ʽ���eK�"�_{-�,ZI����z��[͇�.�̸�BU�5Xr��f`�:�w�IF_�%����|�.�g��� ��Y1������HA���AP��1��+rSu^�}6�ϑ��z�`��?�N�98�E غ�2y����ז7b�g�Ė�"��1�#W9rt��m�J��
�})�7�2j�P:�l�~OR��2wZE���u�:��a�+�S$�>�Đ��h��XS��ʿd�$�+�W�ut�l儿ʵ�f�Y��\$�:��wಝ���`J~��)h�T/59b��T4U)c��OUPiv�M��b���H��U�NG4�m=S��k�����c����Q �0~ޟ�ү+7�.]4CY�ER������w:���ZV4�ݠ����,��|M+�쀚�C�l�K��kfE����|uZӞ�L��`��5U2���L*-;���@����X!���:���1c��K�SJ��&�qƙN=�?;���h�}�f��� a]�C�F�'�Є���XA�k�"�PU��;P�O~KHA֓]s���s��ɢN�Mh�?ŭ#�z��G���v'�)��ʃ,7��<o[��r�/��Z�F.[=%\�xs	�}/U�o��⣺��R�_}�cBC��O�\�w�LE������jt��Ǿ��HtY��k���8��3ЉZ*�n�=��#[L��{G/��ȯ��������P�R�YraG�f�.����w���54����.I��~J�ښ&�]+�!�2ǜ}˟��D��:�^}U�~�$�\����3}�3�0oqMy���� ��p�6k��y������$��e�Hl,M4�d�=�*��(,/�������+���i�F ��S��>�v�rv�$���rw๋���H%LY}�P��̰��Tg��i����_Q�+��6��ђd�r���@�~�XHV�z��c­U��P�e��}���$�����vW��<���X��D�`t������3���8�r����������#�b�C<�%�ߎv���V�Y/i/Y��J�5�g����SW��f���	 >�3��.�a��l=A���u�@�6� q��wŊ���dI
���vB�z�k׏^`�T'�<5�<�ܕ�:�?��ِ�ͫ��KO$<7��0�T���Q^;�p�����}# ��]A���A���Ӈ��,��v��h�T ���Qe-��Z�Ƚu��ލ���{}z4�Ԃի:��}jP&��5d�?2(jj�E�"1��i���;����.������`+���w94l�$�E��u��b�t翤M�����~�h��-VL�^½Ҍw�����"i��o8�2E0#���}^��ŵ��2���?��S��+���7.9�d�����x�V�"ִ��%`b���iA���_��/�eP�t̋m:��� ��&�o�+�	���QY3����o�����]C6D�A�?�_�hΝR"�l��
�:^bUq�C>>�%>mRi����!������u�%d�^csBX����k	�vP��1�M�/�8%��҃��c�bv�-���$=���ݑC���|�k.��xᗌ3�,(�:#�U@Ăm>w �0��a�I�X�`;�;���B�~]���N�/V����eN�g;���Ӊ:dU�{w�A�+�b�C?O��	���`�_׍/�L��<�G� �����*�᡻~f�z6ת9W��R����$�u�j�lo�e$v\tK���񣅌��]���d��Zl�i��`7Ğ���M�9��b�J>��*�?��ԡ����U:�V�9�Mt'�+d��\�,�r^;��i��dt��1X�I{������*Q zܥ����tO���~I�G�W(*yG`w�[�F�S8�ҚP�����L?IJ(2l��{sU���x�f� ��'�� u"9��΃�u�h�7#��_[��]�{�p�'^��GNm� Z�SJ��I]��Z#�5��3�I��5������K��O�0^�"'�-RY[��ڏ4H	�c��tX\(��4�J�s������Ň�KN��Æk�����Á���h�e>1u20�4 �+;!�jU<+�-�1�e�CN�����`�:r�;#������Y̓W�U���.T/�b��6�۵d+�]�,`)�|%E�Ɠ�t������I\
mCc�NS�}��b��m�����ݧ���a �{��P��{(�]�Bf�֥7��*�Gت�N��uP��+h��̏ʭ��i2f��Ė�C_�,y������+���o	�Y�r��X��vc\�H���ǰ��M��tR�[���������3Re�D���x��F���ߜ� ;:�{�S!� c�B�3u$���(Fp 	�0�8)e�?P�}P���f$�= %�����J�������{-r!BH��Q'q'�m����A,��>
߆�ǅ�	�y��Xھ�\^�-�WY�![;��5���s��n��5OfA#��L�I&+�7��Vd�J�+bZ-���-�(�a�y���4��\�,����o�0�	��n�)x �8buѯ2�H�D�w{��>(�?�#ҍ���u��C�׾y�p��7�Ou�-���A�dy���Q������4�v
eI\0_�.����K�"k�m��>�R�]{�p�M�Ma5�2|��8���ě��9pD�xu�}5�w����4��Y�k��eI��f�N�ԵOۏ9�����[�me��k���E�TO~
}q�(��K�e;�u��>+����D��.�gq�?և�b'0�r?��3n��'2���)�#����}��!��r������2���C� �w!.�H���s}�/3x|�9�kb�ˊ(~V֗Ւo������m����(�DQԲA��'�'j���S�����="BDÓ�8
� c'�����
�*����������5��FS4&����hvEW���sv�'���O.��H�-����,u5#v�����M���Mf�X��Ĩ+0��(������X�O�^��m���,�e�vl���/���<�%խ���(�Y�|ދi�d���(9������d�,����ְɰ���mvxb�+�&1���0�ñ�j��7��A����	_�o���X��p$Bz�vP�-�,��"��:C[p���J<,���X6Ny:�����ѷ
�1"�; ���!������"���x�2���&�޺x�~i�2>�	a��d��3�S%
hn�pֆ��~�Y0�]���Z��Kx�wz>o%d�B�&��1b�X c�>���r��ѝՎ��L�(È$�� �Q�f�i_�����_"���3S'�N�3�,�KO���u-�1��UM��_��	���	˘{\TAu��?���p�|Ap �9[L�u�z� �V���l�CC����A>���aiGc���A9�&&Vi��R6�?��K���X�֤f]�T�Z�'R�'��ǉ�\�.օI0��hz(iϊR2VP��-Z�O�I��L�ɫl�kiu1l?M~0h�jZ8�g��q�m��דDaX����7��W��@� ?ș	�����)? .��c�vS�r1ڹ�Fg��w?6�f8�7r�!�Wfn�06���r"���?`�-\����f ) wN�w:(�'��5ǯ�?��!<�K��P���� �`��	����3jpd`� +��/�^K��Q�+�30�Ŝ�iH�\�1�U:TTC�C/�U����ݎ��eA)��n�tbZPU��{���B����bp�O��<.S9��$qڴ9���r$v�G@qˉ��5���g�j��5d��2=��7�*D{r ՟%f�(`�@;�B2���Z��;���UW�[�xԢ�N2�=ꕤJV�Jg�����a�!U����)�4'j�?"�iz�u5tM�� hV�*����@��#�����W9��s�0��J��n�b!4��_h����f>x�V#��N�_�~����>����Q�dqD+g�9): ��dͿ���ơ�DH�"��ax��Ra��;�@�|(��,���1'�!7O�|��v���y1+ڸ]971�1���9�Ee�HX~��7�3S��3����y)u�����C;�rsQ$��Ў+��S�D�/0�t+���$6j���yN���B��Uϔ��N�0����S]R�VS�gq1I�Î9F<�i�v��Y��2D�Qֶ��P�S�Tی�9q{imn�:d��A��W~�p��9�`�+h��s$7	�A�D�{lR�-ϐ��h<�|=��U�ٖʈ<����� V�d2�W����g��T2Ja��}o���=��_���WiQ��*I��N ��b��U�k���X&�#|O�<e�?�h!l'ݿ��zg6��vE��!��!�:8����ǇqD���A�Zs\���A�hNC���|{��{ N��0r뤠s��l}������	_s��3��p���!�[o��:�[$�,�'��3�v)Pyj�U�W� hc<���߻l�j#���JJ��wV���K��z����J��+[�	���Bd�t��*8���Z���� �09���#��#{p�Z;$���!�^
SgZ�X�Wt��l�r��+V������U�I��¸"E镸���ҷf�s�i�W~F��U�K���nl�ِ;�vw%��T|�n�B1�;�����n��3��00�Fpf�A����r^�9�,�œg$��')v��v��X���{M1��M�l^�4(��y�g5Ъ�`�����?\ݰ0:Q����L�D�{�T���X��>F.ϝcN��F��+	��Zl�,��A��wd>��u��A��a�PȺ_eX���UaS$���g̥�_;n��]!b�5T��9�����v&�9r��;p����H�װ�K�uR�sJ���.;\I�=��S���s])�O�|��^�cvO���NGe]���
E��d�뿒��A����N^F`
�ך+����TI4��Zt���op�!t��#�����!
}�?����X�e���"
A�V�:i�E�o��)��ҧ���hq�5�쓝�6���M��Q�̓�:����3Z
��ؑN�t��o�ݢ{@:�|,�!*\*�9	)�
Z�H����q����h퐩h�hW������a�?����Ľ� ��TBv��s�'o�GV-�OL�	�\�䴢������l��P�4p����7y3�B��$�;O�{�:n���M�]�5�Ĭj���gͺ�r�aT1mL�6g��e:��+哣W`C9�؜�vx�XV-�!F�A�i#æ~��#M���#�rlEL"��D	z���v\�
k����]��u�sء�U�<e�W.�W@�R1v[�-� ��˵�0wt:�T�⨊�4�O�*���t���SVY_~Zx)���7N�*0m�䙨�:p��n����!�Uu'℟(�|g!-� �L/���F�AU��$BN�"HNo�phY����X�ƻf��b5\�+F�n ߏU� vl����2�_s�Y�e�j�5���n� ��N���a�
ֻ��LjZL?1+=}�~���VQ��Y@�hd���H7H�˗��cp�RvB�2�����25�rƸ�z9vX;C95�Ѡ�WW�q�ă��X��=]nèM��i��
�Bbm�R��0�O���C�l���	�s�=�`�^�0�^&D�^��4%����W�'�sB�d,������V5'�ʆMpR�u��@�
/�D@[���9����˽$�[$W��y�pZ�QW.�� ���(���#Fr�;�v��9`8�4��`"�z��9�5.0�ŭ��4�ް�9��e0��������h��7e^�F9gcF6��h��)(��@�"إ��qē����ұ�mnT4�0�vMxeŌ�뫅=F����G)���� ^����O��K����TAb����J�6H�ي��C$Pw1��[e�##�ɼ�9eҍ���`o<�D�Ѯ�{^����Fj�t��=F�������_ǹ�v���幝�!A I�	4��׈5���X<��h@X$��4
��_��n��\����o��F�n��M�ID@���-��XS4�����F9���us��:(T^m�@khY��{8�<@A�nޥ�Il����Pj�uxMb<�M�)���;�A�ͧ�>�z���m1fՓYO��j�x����E��]�5�.E��ySrV,��8�ֳD�P|��Kح=e�	���S!N'�>��U���C�=v�A5S6D���� 9ɫp�0�=�NՀ)���V�e�:u �eu/vI����mS5�]>�A���4�R*���

�Y��zSЮ*I���J����G3��r��G7�ig'��!m�T#��ғ����]���tO#�Y�{@�P�1N>��݈FK