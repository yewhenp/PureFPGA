��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��㙂��c���љAtC�~�<ۼ���U�"�D��([z>��(gR�#���Zf�J�[���OE�X�#����z�3��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ�Goo�27Mӗ7��� 1!8��,/�RV�6b���jtTEfm=5G��$�������M\�w���ua���0aޮ�`� /�x.�Z-ȮĤ��� [b	�$��#�n�L�Yw�3Q�g��a0�ܜ��ū�1�Lߪ��v&ۛb(��[�]�j���`�.AؿU9#��F��<�@v�$��7r�B��0ؤ�2	��	�Y�{f�����^�LY���eCMG(��P�&_�Y�^���{����T�K�W�"r@�������Z}yrq)Yٹ�����>�_!���tm3��{�E�C7���b2�[m�����A� �$�5�ڬa�8�!�1"�:�4G{��	���k��������#!�c�GڝYUľ>�X��T�p]�T�R�{G�U0+E}��'ٰP��Q�iK-���d�ʬ?�m��9S�v���m��rP?��n4֣�.�k���w�͆�{\Ф���1r}e��4պW��"׎7��͛(�(qP��n��.CpP�)\�����9�Q����M���mI�c3�l1Nq&���Ht��'ȕU�,O�f{�%=
\�yJ�G��5�R�l����u���'�6y𠹗W�s@��ʿ^|O�7W��@'�]qD���X@�s�Ud�]P�g��]K�5��+��i3�82!���p,���a�U��>A�J�U�)�A2%Bz��y��@tx�GS�|!rm���q�">&g'v����m@I�̠�, ���~��6���IF�ɢJ��؃p���(t��jN�������� �ܖv���7_���H5!٥9��{���J�����ԏ�|B�췰�Nzt�Snz��b� �@�EL�)Sĩ�y��+R��ޞ0U��U)����ᬘc�zw�1kCFR�� �:�C2[����<݀��#�����j�/:fȪ5/D�������k[�a
Ѓ'B�IK�^��s�j쒬��5}xS�0C����2u�_ �3D��6޺��v�wBZ�U����n�� �7SӅ���)/��g�_���N�f*Ų��,^Q�rb�\��DKVv\��&�W�F�C�&K$���?�v�~%"�g��̆uh)�oN�咉w@�7H!�F��H��g-���<�f��1$nJ0JSg�Y�i#f G׍�*wp��)'tt�� ��Ԋ����8
	���aYI�)G60D1�o��q��X�F�?-�I%�؇'�"}w>ʵ[��۽l&���3���d�۷�I��D.M�6^��ku��朚���r��6�͹vy��/Z�8{yI�w+r�y�[���,|����1K&T��G�4a��R9�Z����_>(�w���I��S=	/	(��*\��� �c����!�Hf�p$��&��|��T����a�O�}����C����j�Iڀ�dsn��<Ppcc;C�Ad�8Sw���5��r29%��l��&֦<)	\'�Ɨ�3�aͰ�Rr�֯���[����y�t��K���������I�5��=���'����`f� #�
��{����'�·�\��tr��@�}��k-�b5��1��B���oP!;�U��\T����1�꼙WU�������?�֤E��TJ��.s��D�It3�FS첞h�}��� ����������*dK��o�������j�c'5�|��๿�t�"r���"]*�7���Q����� ��tF�8��t������}.�h�\�'�P�5�J{��o�DX�%�
��_���H��K�B2B�Q\ʘV!��"oq�|�~W�rА.9qK�t�q���@�,R,�h�\�~b� ��n��G��܂�	6�k��8)�� e��m`WȈ���͇±��&��fҀ�
��y��B�F�t8�N���W�p,�_��/]�L���������S	i�,@��]�1B���,]y���)rE� �k�j�^q�=��=r_�2�ٔdf�*eF�__�S�3�t0���ߤ�7���Xr���� ��[F&�I�VtA*k���0�{$n� �9�tA��ӌ���\c�_��B�
�j��pX�5d:@�j�{�Ip�v�R.b4{>j�zu.p�0EIϔk�[�ƛM:ڄe���|u��aKe!��*#�r�1�k��nd������QS�#��-��&-�W��6~,�&�M�6f���t~DK�u� ㈺�^��#X��,���L�1d�
5̀��fE��6i���k����)�1o ���X-�'�7Es����7a"�*�'�Y�y�D�=>1
3���'��|-�<ry�z���;>l�y�~oTΊ�<Ż�U%�ЩV MU,5�T_+�`
[*��	�����T܂ ��\�8�V��Q����4�,��Y	(�l��:���x~�P|�4%*�. ��S�� ���Yy}޶��Bdt+���v��b�E|=k�ޒ� .����l��$��8G�h}�u�?d��h����9Y��@(�t��$��F����#=m�v�h,yq�Re�����j��V���QG�)��|>��@$�ӍN7�ݵ
P_0�������zG
��.j����I-ʮ�����v����9�L�$���d��­�z���V;�ӿ^ܰ$���δ�pb�]孏�Ә�蚵W�� �@o;v�����N��ϻQ&s<2W��,UB�N$_��X��
U��
J��)���N�/`�V`Vmг��>�'�,��{�����d�v��_�1�_��oM�DŮo�� ^ʸ�	�od�s�Ńu�;�J�����j��D�s�u�6$����@��"w�i��w��1���������̶�D8���Q+����XЎ�W,m��&H#�YyZ�U���v��w��l�*n1�z��/
i_�9�~�*U�|��Bq���TM׳�8�T�)�T\������EiNOC|D>`�𶻆«x��}��كץ7��G���l�m�s�d����?�!��$
<8v�;��C�Z�/��n	���=ڊ׺��l`5��i���{��>���D��1�OBJzbW�'Z����іV�����6��w/z{�K{��b4��wx��$Y���*���s:�W-=P����Ʒh�r���#hr.���8)xS�I	�D;^$K��jWg���L��t?���>FǇH�2��YZ���$��t�ԣۆ�0o���:��=_=���;x�'?��Pw�qM>R�xO�1��>K�ˏbO���W�;U�6�������!P Z��7�Y�����T��$HU"t�O[��k\
�}�J&plI�Q:�ds7[|��$ӣ)���Rl��%&�9J�9~�=�Ǝ�[�q8�KI$ɉJ�f�.�����¡$�6��Fa8� b�v늳�'���*���4%#��'�v��މsSل�>�D*hg̪ĭ�H�6�$�P��M�XS�}:��QE*���M�b�*�H�A?��^̉R�o=8==�Z�	m�6`����t�g��vG��x#ǫEC#@�X#��⁮�HNls�Q��|N�,��������&���&5�����bAAl���^ܟ���/#<�M�����8���@�
��`����V��9����%��U��Ѥ�jLqT^�����PP٣�'^���0|�E�7��Cb�9o�~�0�
1��]Nn��˔mL�'�Uȏ��L{�[�N$��w��d!�&��X�a�*�֧"+<Q��N3�j!i��-�F���3X�w�l��RGfj"��AA�����5��� ~���#�U����F`e���e��E�b��o=�;��k@�.<~�
D!�*�3����'^@?A�Cs�����g`��z�d��f�C��-����JjaXqt�;����_"�$�k�T���G�9�%4ݴWj���������7�'h�-��ܿ`Y���d|�/[�7��Az�g�����xܔǢ�_{��,�%ۚ��i�����l]�S�[�!:�1�K�޵��@z��9o���,r;�y"�*Nj�c3��O��-j�T��2N~�A2O��ڡ��A�y!S�Gt��'��m`�g�4FSd���b��O*�V?ΚT���8�9����/�o��.U���0(Q[�oF�G����c�yH۲w���ǰ�I�weI1�BH���]T����{B���@;�m �"�|7�����'9�?�c��l����]m�|W�����r̕q����I[I}�,���^�A�Ntu�GFF����Be�.�n�������E���~.2Sɶ
R��7��V�术	f����y�4C�Xh����/ꞹ�v�)�v�^(�3�������b��)�f�@�V�U
�G��d�t��7��Lk�vϗ�G����r�`�