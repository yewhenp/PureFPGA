��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ� �t;l��(Ur�D*��3ad��Lt@�2�.��iۉϯ����I��s�:��|�L a���W����*�w�-kf�8�T����	Gy�-V#kx����JvEW�'*q���順���T.\��eF!*�Xx�1�������r�LL���CJ^�t�"�̫�r�ïs�g��q�/��T�7�o�-W��=j��������z��a|6_x&\W>�XF���z&�ہ���F�6vtثy�n!�0$�	�Y��W`N�!����$l��Z+���R���w��*��F�i��C����ry똩a�GuW�8j�Ս��h����<�˳U�]���-�e Yx'.%ytN��J#2�z���b<f��D��:��43��oUr�1� �|;	�p�P�	�~���aj�I��T@��<�D/�zmL� �,˺$�/��f�0�Hb�JE����𬇯��3���^�Lz���[-5,����O�(�-�Zc9���w?y��K�T(����y�����c�^腠&�B���`^vg���vպ:�F*�L�d8)R���'E�c&L��y�vܪ���ql�m2�I�.�
�U�0!�P���.�lb�Sz���]�7��Og��MPE��A�uX���,�%]6�teiz	�]�3Ë�Q�.�ZFA�>�i������oEv(�&jđ�TX��(��le�H�ϰG�Zu�J�SO	b�u_`Ap�[3U��h݉|���&Clz�?Ŝ9��ڑ=i�GM@�	���x�Γ�aZ��b� 2^?q��>0Mԑʩ��>�����5&��������Z���s�m�tO�C��u����N̫�)-B���Pqvt�&l����z�Q ���$x�z�e@���n4���.�y���ϋ�q��j�/-�w�,�����=��MT��p��c���ԛ���Z�Z̺�r�_��KU�=�R�:`�T�F�3�6`y�}v����s]�42;�"��t��"��x��#��9�=s!�����q7�a��5X0��|���C����;^�bhKm1����Q��o���sn�#Y��;��&�
@��*����w�_=�#�$���8�?b�#�q@�NAҿ�з��r��)����wt� {��ds����X���7��/L���p7�e�o���| �#��ǂ�� E�^���
�k��z���Ǵ�6�p���o�{������CI��`h1��Ә���af�T���B^yZZa�ڸn���w�d��P���Y�\h�^^�}ܜ�5�֕��ׅX�򛃝>��2V��0?���Ɓ8�,�	�>ԅgJ�����M��{v��W�����"�xK���� ��5G���}kӋ�ˠ���]�'*�����5&>�c����,� �@�$�S9
KjsS�	s�2�U�)�^_�k;�P%g�*�OS-x�ԏZR�c��/Ä]�'"�/`���&%���;�����9�+)fr��|Ih`���yT��Fl�p�yV�'��.M�#q�-���]%(�	�Ún��^��LLax���%T	8MP�Z�=c���J
 �t=���I)K��::�����ᐞL|�	-���/!��أ2ޭ�j�O:O������g%%�����ش���ѩ_�o'��9��3�!��.��������>cPT�����S"pzY�8Q���i�G���$>ς���
y�DV_s���V��8
�F���I���������Í�E?�g�� 3E&�~��v�5G��Vw'� /���4J�LZ�0^��ܰ�����U��@�]®{O���G�J�6��m
�����`-V�o��6h/����M��҆�i�R2�~�1������!�&x�!P����?`��gT����x ��!�K��E���j6̅������86%"!�H�OB�1�rZt<6в3�%�͕!�Xq�T�BZ-���)M&ɚ������`5���w6<irv�O����N��ۙZ�e�!��Yۄg�zv[�t�n��%��`�v���6�݋k~���@N����;YB_u{��SG��5M�6���s�%��]7�6a�q�(�D�����~[|���7�	�(kv¢gW��f<�<��6s.ʀ�{��r��60~�r}ñ�L������e���R��T�k��/@	��L5�����wA���Ok�Č��e�۴v7�E��E�p���f��C�"���S�D��y	��� _?�V�Y�S4nU���ݲ�`$�ZB`���O��4�Ϧ�RE�_��q��/����fiz����O�J̶���
̉��.��Q{)3׼���%�>/� A�@����V{�|:f*ڈw�1��WS�L�{��<�6�	��]�����u�V�H7�
)嬯��+���S�b��H�V�����g��td�//�u6ڧG�#��oU����V���VM��̮�|H�,N��L��C�q�-���
,z�?�����6Y�J|RA~�}���5�y�`[u���Qw�1K�C.?V�����It��T�VY��۔���t�������$���oWI�tCCκ`V��lG/yt�.]�~�Ul�0!���W�{�ꥏ��u��t�
%�/_ Z�hB���4�.;�%,�19�9�X�oz�,�G�^|<{�.1��M(�����լA,�U5[����;:����Y�+����Ƨ:q����l4��iHk`3��%d	�����S�곢hmYɃ�o	jn0�'����>ߵ��������P�l�b��2������Q��H���C���.�� �5�=�~����0v+�|R#}4Z�-�s�����Q�A)n�d̅������az%��R�T�J��x��%���>�~q<^'���e��V�&�{m�)����d�q�/��F��E�aG�+\��+ �����T�Tw㬀S_�?k�L@�~pN�o0�N���o 6yrȅPȽN1��-��Ɯ�)rV;_�g�r�4�~���A��鶹!��L1;�J#��I#������s��p��i
]��Cy�9���'Q,MXիCVĆ��w��a*�*�s�a Ǳ�b��w�����4��(D��p~(�$=w�٭�y5W�Q�!lB@�O�@��K����]������R�����!����o�k���d�v[	�<�y�U�mJY'�ـs�*o�H�e�a��^Pl�A��RO�W�[��&4��o�/?�u~M��`T���_;�>�(gmL)7���-1�k_P�RH}�Kj��Ha�tx�6g{�L�ѽ��&3�lc���YDA)���^&y	�h� Q�&�ޮĻ����ֳֻ�u���j3��]b8Y�p�N���c���Ϻ�6�+pD����K4��Gcaq���L^.<*8J]N�&�Z"q��|ޙ�`N9�S(��Bq(��;x�!M���ey��d/|`�.��~����$t\�����XW�G����s�AN$�c�;bI����A5����fҊf?m \�ى���m���"V)8�PI�4i�Q{#�O���IY��F{��Y��$���W^����k��ҏ���Mc?�I����#E��*��[�
k]def����.N��jG�
s�p��dW����I��يx2\	m��K�d#�2R�V�Y�Z��OfJ6��Ì���-��I�%�T�g).�:�`����JH��-�7^�ˤ�Ƹ@>�4�jb����Ec]zb�q$��e/(Hf|��3��&��\e��K�H��F���^2���.�-�ȟ�7s����;��
nZ-�9�� �B
d)~�ʨ(#Ee�t)��O�-�BKE����Hhr��|ٗ8�%��#��V��Q\��vD��j�c���(��e8�N,M�� ���'�&�#��r����v!��y��������Ch|�e%~��t�8;������C~K�MI9��"
u�mH���[7$y�Fkޙ��V~��o��z	���>6T����5�tk�I��k<ϙu{���>ʘCs�k����su߼�[%.k2G�8= ��3�P8�)�#J�6b��S%#6���Z�e�Ňs&��:�r(���`~@o<s�I�$��q�����gyp�69�!�=�h�a,L����ZL{�M�A�C$��	eN��X�J��܌�_��rϛ��6_q,�ڒ�6�<��xO��BOI�mMW��h?`�Ɛ��A~E��{�R�K]���!"�r�9ʪll�Bn�o A�g6u;$lIᣒ%{C��>�|�5��KІ����K(�*��?\^ࡵl7Y�������M�qg��t�3Ġ�J�D;���v+�2&f)w����v��������1�����wʰ�־��������9���z
�r"�{�����D� �XXc��?CG�����q5Y���6�*3{t���Y�}ewVy.��Q9���$����a�e80դ�N=^����� e?~A�s���94�|���?�Ǻ)@5�5�axoײa�z�0���L\
�zW�6٫��kz&n �}3?iCjoU���^@ѥ�ߩ|���he�䇹�^�k�tĽ6Jc�3�5�I{��b��=�j�܎l�#ʅ,��d�����#VF�Ӽlú>Nh���Nu��	��v�c�)+�KLǭ+V����%���9�݂2J��/V��K�I&6���G�����1twQԺ�g7�3���0vۉg�YoJw��Vs�����o��%Z�BB�b�D���fz=��8k�����a��j��gm�2�����"*���z������Rs�8c���2���G��[ߛm�4�����NClߎ�"���[c��W�%"�.\e��F�G��V��*ԯ������Mu;Z\�e�sV�?e/�7cH`�!��o�����;#��[�T�C����~N�q�9|�������z �3����*>{����zduU��:;]�`���B�C�fC�Ś�?ե49��(	�͎)Җ�#*Y`�R����KK�5�+H��<�0����X=]~uϪ�{�a��2�?�X�Y��tR��TX�K��4m�X�e2�(���KP�W�~9�p�ct�.�R�O�/b��d�ϸQ���~��xݠ�!��~���>ҕ^{���| ����	;���p��n?���4}+��<����vԕ �ͶY�_]���]��D̛o��3(���ӋPB�y����W�$��@��L�f��e��JS�!<�]������-{O�r]9���㺹v�ڒ���k�u��}�Ȥl�I��Q�Ќ4V�a���[�������ԝ|k,e
8�uE������E W�*�5r���3y�p`zo�٢�<͇�D���RV�LJ����@�����N] :2xs�;��e��/�i������,�4�?f(�������C"-����?ڶ�d�s��;m�f�N!�+�塴h�"0�Y�Vl9&����b��
�I���Wf��_���FL<�w5��CQ���O��D=�M.ϡ7 ��l���q����7cQ*xK���.ww�����@/Nat�$	�����<���N��g֔&w%�G���KD�L.R45G�%}C�H
��;����������=y��,.�+訒�r/��P���?��ָ�lha�
q��k��z��t�۩@isO�y$�)#�����ֺorU��^�?��ۜ���4�����c�f�]�qο��S4�|'�u����$(�!��_̮Rm;�)��u�G�����:l�g�Y�e�[�"�Rq uþ�ﶫ>�O೾�'�(~�t�^⟔����.@�u$D�݋\�hJ��1�O8m�ϩ1(R�/}L��=+������W

�[d�C�Z�u��$�:q"����}%��{���Q�#X?y�5�z�%�Wp|��o�jb�cW�L����H� 8(�F:{a����>k�F�Ttk�|L~������E���O��Y��5J8��~�2��}��Q�z�lTQb�/ W�qQ��̮�rh;��l���pG�7����-A8��RƧE��e�7�NC�!q��'?ı�P�P޴kz����� �!^!��#9%�f�9UXYZ�Ԁ`��!?�]$��~e�"���!�R�͜�����q�q�s�Ӣ�h���p�'�a�#����5��eq�;�u����kI=m�`
���^f���'�ߡ����M���EHUt�Z�����hU�/������6@9͟l����&u0��A#Ds�˝)	�5����$f_]���1��Ḱze�������Y�6�h���?G�QT8\�'w5^�&��FB⊖����zC5�c�!�q�?�u��_9���֮n)j(w�z�*������[�RTY9H WԔ�>/p2���u���UR�[Y���%��E�|�����0�?�)�+����~�d�7aE*���L������_#�yؗ��U
�����Z�:2��=�K�����(#8���v��Q�3�i䂵���C�FXI�l 6��� 6���z�h�[�Q�z��|9AMu%���Kx݇�B�+(=&��h6]�Im��rX�G�g�f�C=7v���Z����;ہ��Bܡ��(@캟��!ZSg;��)]"!cŶ���fo�"L�X������)^FY�����&d�+bi�b3���x����%����Ƴ<'�B����3"N�>I��:m��1S���E��'����Ċfoe��E���F�n�>>��r�ݦ�u�[xC��~$�s�����k�7AsG������aX�JG�� 9�\���(`��h�3�jU��G�3]��{��Y��!�p`7G�����\����r��������,w��T_y%�Kф��cS���)6ne��x�)��(��.ui��������x#���r�y\�ڮ���2�Z��4�-� I��-x���{w�ӣ��xH��Dar��_\����˷�&r��l֡��2?�R��ɽ����fls��IN��31R���,i��ϩ�'�Մqw��7tD�w��]����V�rt�H��Ba���"��p�~�6��/�C�ρ�����,�tmZ�M_ +����^	�䖳� �3�P&�t���J�:y��L�YI��Ɲ�#lO!_���I 9+BVNNd�[_�{r#���c�=���u�^��;2�D��� �F��~�2��MЦܖ�cZȚ�5O(>^�d"w���Xfm[�$1�S��)0�_�f�r��?�*�a�Dl�_S��������F�(�j3�V�I�՟a��jMzwdcA�x��@m���Q���oA����ݏ�i^�Ҵ����p�|p�����x���r2�ap>zz��g���2%"����$]^��σU��}��<}��3�t|��*U�{�QȮ��8I�'��!�֎����K �Cc�M�1Z���>-%�h�d�)����)O�����$��7���5J)�gf����yt�%�J�*!�0�X�y�_z+r!@c�T�u���9�<��H��T��Y��֍F�̭j��ժ�H��M���*�z7P��s	{��U��י��YW
����.>u���F�"���l�cֿh��!W�x_��Ёk%A�7w���'��ew��o �:a V�U���:�^9���'߯#��3ߋ#^x0e�Y�� d�YO>�j��_*��MQc�T@-��l�I>:�(ʿ�	/���@������r�^O�u������~�Сh��Q�����'���)����vM�a8����ŹfKЊs�Qf����GVӻTv�I5�?���" ���� R 9������7q������;g5��O��࿫�9up�d��g�V�15�d�'j1�4*�3��|��nM�d�� @Dy�
j'����y1�O��/QU0�uwnvk	�-6�F>9�R[��?fv��G��Ds��7��QS�o���ct�����/?G��Q�~RĨ����`��[��ݳ�9uU������x����@X��Ov%�*7��k����ͩ~�E��VQl4�cK��N��8Ҕ��<�Et�*Ƙ�̚^T�Bgl���w����������x�@�9�R+R�$m$�����J��!��\����{Q�Fx}����$j�������"�pזh���WF|����~K����
��eע'�L{8|Q���b,I����Z�ұ��+vU��m��Q�F��}� �K�I� f�?�E-��6޷�"Xp?����(i�Fɵ�ҧ�k���Ok��?#����g;��$ȅN�+�LX�w������Ǭic�i��R�n�\���Ι \��m.���8!]7�E��D�&F_m�����L�P������/s���Q��a+�WĸaI�Յ@���L���1s;�;И �:F�;��W��b���I�|��.�;W9��aW��Fҷ���IG�ٞ�)e�)�=�ĩT�<�Xf쎟�#�ޯ�M%���l!�oCv;Ɓ#�����)�3�D�I�
@����}�2WD�������,�Kјj)��Rᠬ$��������j3��9�I	S��al�� ^�B�j槳�Ʋ}J1%�L|��Jr��R��ӧ�w�n�pٯ�/{-S/����`�U�$p���I�D����VQ�T]�7٭�d�ָ!���l,q�L�5���l௟�m�����'���H���SH*�룂�ɜ�������:)bc��i�dM%��Oe/9�]�h���-�>J���߹n�����0�����1�k��%ŀ���%�m"�*Bn�d��h��z5�lP,���4�|��?����h�q�bT�I������a��G���F�c�3v�e���P1P��� ����WY�n!���B�7���ǦV�!���B�QR,���O�xk:�_�i&7"�;�w�d������1��O��
�S�B����Og]"ش�2�ws��-��\15������{9�i~u��7��k&,%#}7�0�x���a��j��-�Y�Y��lu��{��KQ-����`2���v����T�B�ˠ��yFd��Y�q�j8p7M��
i��T
键xGc���8sr�]o���r R-Y��+�~�	��lJ|�����!��x���%�������+{�ni ���2j��u���Y���|�����;&��MԐV\�����#g*ީ�몄X6]���hc~k.�6�t�5E*���=s���y����5�~g��כ8r�� !�+��B;�{t6>�i}��uo�gl�/�Jb-���E/n��g�y'��Iv;�SD�-�1J��`y�SN�]��c[8��	��T�$|�
ғ��I/k{Y'لk~�.� m���� ;Z�[��9�[�����e�������=  r��]N
\F$"� ��yA5��H+��}N�,��zl��O�8�;נ��3�s�8��a�o?��qO��x*e~䣈6��5~����ui�j�v`DYM	����9��^	N�Y�K%G(��5����"���KZ�8��5�������Ƒ�k��H�${�GR�XU1��
�a�K���ydь��9����֋Cz��PGr{U)�Y4��1<���Ǳ������㊨�$r9Iؚf��ӯb6�@q��%6�z?a��n��4��p�B5�I��-���#!�,N�'�J]_rG��>)�Y���k��Y5G�7����91�j�K�p�N���f�S�s߭<�y�_\�����r���j�p�&�����KqK<�jN���{nv�7���SR�0DX��zp��M�
�)���½',|*]!�?`2�l��Q⏱8�h��R=�o��S()$OW� ���$N�5���iRɛ5_ �� Z�(�%l"��f�E�����L�JoC��^���~�)
Hl ��'I���#��|/�y͑%�5(d�>�Zd�7%r-VO�cÓ�hҤ?6��6)C'��. �1�H9�Q����#������_>�
�9$�{�ʗ� [(W�g���s���vG��0ԆOő��G���"�e����|�a��܊<���T �7��Iu$v��q(��ӫ�D�G. 4 ���얷�z� ���U�
��Xm�#�i�j#��Uw}�i���6V�Ҧ��Ȝr�y��f�q\�hJV�SAz��ޑ�uG#ʠ*\����F���+��{�tE���y�����<��[㝵�����I�b1#V���m)�^�����gON��@8�}��l�f϶��1)>'�#��k��w�깠�s��-a ��:R�[�jm^wQ=>&���pU=�9g6�����/�y�lm��T͍��r�bgsIT�����ythիtQc%��4���S<⇆�S����r����+���̭S�*�`;\�N�(Un�S6a� ^��M��7��=棲!a�F>���n��/(#�>�=<9k�g��#��s��V#�A/W2�������C5���]d��J��~c