��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_����]ׇ5�F$�,M�6��"�����hgu��:?)�V"*�T��2�6�v8,��Q�3"S�Ƀ���+3ӊ�ɽa�xw�W&���K(�j�G��O���"5�@wu��Yq��ٖ�v�k�K�\p�	��'ңt�>��qRޅ��/r������Cu���Q��V�+��p�A��WAV��O� ,ӿ�b�Fl��`ǔ<�~�ىs�@�0�%21c�*���(V�V����IG�7f�;`�
�˗x(n�0��"�%y~��Z�� L�o�D�y��Nl������W��/���F�D.1V/%�?��J5�s�������t�zDx4�@�V����鞖�z뻣Hڢ��1�b����3�枓��X
"��e����o����v�6�Zy��sgG@�F���9c�B)��7�}�x7o�=�G�� ��=p�r"A
�o�љ�u��C�aߗ��a����I˚FB+�<2����;l�}�R�9#�n��#	�dE��UB^^x�����4ʵ:STcF��M?*Jh��܊����e3~���yYG��f
���Bh�)14e]�ꎧp"�%O�����J��҄�kS��:��gܱa){�n^t�(���Ձ��^Qo|�����Ā>�^��7�n$�	r/���4��Df�Wkjy�y���V<���ڬ���Y���@Q���z�d2���m;TT�!O����P��]��2{��gS�w�����J1-?��v�u&1s;D�l�\PV�~�X�3Y���	� �٭�뙬X��bܱ��2��s�����*kll(��}tO���iO�� �b�*��.2�N� Y����Β��e��@�R�^��(����Eu����6Lg��|�D0~���r3��0N���|٧ǂ�;
��"+������`Y�Ƴ��E�ϧ!��#7i_�����&TȼN�F��+�h��/nn�Nni�_]���P`��+XاS�7���&|L�-��+�3�(�b�Vz���� ��ƩUnD��<C>7Ĺ���D�Q1A��,ե�;[�x�B��58/�C��a�	�?�H�������9�m���^�A��=��Ud�+���9">ۏU-/ˏ�q�R�/,}9�}虴��9�@{T�O�o��u[����T��C��6���,ٯJ��Th��t����n��e�\W7�T"]Ȝ�w>���kk�;ʹ��ʊ`��\i�3\;������j�Z�y'u�KH�7�����<�[�[�>C�b�`f���a��G���Ĵ�=���J�O6�*3.��S_�f;޼]0�_��ϮF�IU�<P/���y�w5�"��:�L�r�p��%κ�d�������a`VȌ@U2�[�����T��j��Z��X�h���]�r{!T�]A(�p��Ǆ�h<X|�t{�3��C�?����J�^q�v���_��w�U���{K7p��D��$���-�Ai֝j������T��U?�)�~�Zx�kg�� ;��j2Cz���L���,B�A�GS���mb��fd��Y�Y$�	!!�fX3�1|,@yY�b�vM���P�K��x��UU�2���b!:��'	���OAL������י:��@�1Y��c����ZL�k.��"2+��e�4E�o�py��$��"Y���M��&�������/�c���:�:?�,�_sbqU/,�{�z�`=&�bH�"���C���K������K�usd���[ɹeR@��j)?�%�"�~����e�"��-?�;D_Ä�_rTSO��-{�����o4���_�簦���.Ei�\����ʠ��}j� %�x�q������!vFũ��$�m�$���\���F���;&�~��͊�jbt��Fݳ��aL�fr|5�s�i������]z=��e@�")����7���d|XݡaI��b��.T���������>>_���&h�! �u=t*Od-��k9&����A�z�S=7:�)L�`��7V��2?v�L&XFY��l�ӿ�k/� c�w�"+��)R��ӗ�ߙAx!��(�y�[��R1W�Dx$o|5�.z��f޽AA~��F�G�X�ax��B��r"�f�����/�{qĒ�u\�q��	��pqw�Q�a��[E ���Gڦ�B���=��S����l��r��㑁����X&`���dR	k{v=��m�#Lzx�e�,!�k�a��/3MWC��/�e�9}�����eAY���9��D[̛ ֠޻Oݭcg�"
D�F*��r�G%�
0�_xK��f������L�~�Ӡ�r�*����A�taS�I���:��jqfw"=9�%���+��-\�.v�#��E��g�V��[>�W�cT������a�7�w��
;��x������ �þ��F��$v���P�ǘ($�n|#9S���Z�s`��>[
����w5ߴ2��Jruƃ����#j��r���p+��Ц!+
�"���P_�=�5H"j'�"SL�7D�N��G&���S��.Y������%�����QC�y,75W���YR��6����h�Ϙթ�{皻�]���>�ϧ/�0�ƣU���B��M��V]��*���^�M�)o2�"$��D��H�l:k�����������S퍮�6�u�=Ĝ>/�-�~��kDJT�z�ω�;A�Qk�:D�5���P���-��Yi[���c��b�7�^����V����o���G�3g;@Y�	��*�3�Ѽ3P�շ˚ʱ�4�[SY����������8�b�D%b*�5~e����IS �Jђ��(��-b�D�2��V���%�w��)_�ن�+5g�E��%�B0z���s6@�J�K#���/����̶��E$Э�����Vk@�u%Z�5az1�FV�^�a����5P���92�j-\�������{Ϳǆw�ɺ�_:GJ����e?O�,�y��j�Лyb�K��)�s?Gf).$Z��*�?L��#Nt���G`?|�#P\���:���D_�x��:�I����4��7۶��L�6�^��	y����}������
%3��}"��fRϼ���<x;��/Yv��,���V{�l��O&d�B�]ձ1��p86Q����P��>)��hZ�1T���I���2�Qf	��)��X���w�>h�WeO���;N������þ��f��	�����$)Y>�~�ʱ�e�J�.3*��S������\�L[�<AF��Y���ܝjZF��O��\t+����;0�4�he	l��`���]��t`a��SY�.�.L�c6�=Qz]h�PIU0�[�dO�R�nbf�ӡ��u&��<��t�خ��������� UR�=I=9v�cL��o�*L�K�'[b�#�jt^��5}j!���82�̳נ�[X��(��3���|�?a=���Jo��B��hr�ha|���x�NDgdbdp(��Wvݶ�VZ��l�"�PS�ǅl�F���'n�ޮ����P�f��rh��y�!��X�)��Ux@�2�Z8��~���8+�dh�8�Y�np��~B�η���P_����W<�+�z���"��
�*
y�1s�f�g�߀<F�U���E��X���%<BIʹ�x��en���OW�:�iu|����5}�[F����%�T�(3ċ@�u@+"�I�t^��#(O���.�nZu�X|A���̮�1&���O%�[_����=߂d'�&¬�)d��D�����Q׉��P�G�E�\"b����T2�7�J��B�:�*
�L���l��uU�Q��1��ywK�_ �爉�ʂo����CiPΩ.���Xo�\�UH@E�1��>�F�2a�ي��<�~^hOz�~�/�:G��f��%�В��.d�V��{x��e'��!n��.�&J�|T�P.��$�'h||Z�Dp6n��p�)���
f*L:!�ʟ_�m1����p^b@L}B]�K���LH,� 1��H�����+10��nא:e��C�C�}�]��Iɤ,?VZ ��SԔ��R�E%T5,x�����4��B�cG�T�-�;5�N�-������0K�Q����+�yK^�+���%�{��$Š���\.��w<��'0B�����&��W����S>+��Ӕ��f	ʼ�0�@�;�Zh�鉁?��_h�L2?3]��DD_�bcJT��o��]���ќu%Mɫ�s�4%mYs|�����*s��9�;�)�j�lG�m�K�WDF>�����f�~���W6�>�m���t�N�E=���JњU�����^�,�R*�%_��6��X��3�@
a@�a��ѐ���,Bq�d�{8�lF�4F�-�
=�^����%��B�����A�����׆�5(�ǉ�$�^>1���b32j�qEEg��N��`���؈��zI���a!�H�,��U�kr�yw�8Z�	I���M*��R�CX����]��
�7�k�Q��J�B��S�,�@Q`kѰ9I���^�p���·��GU�V��+4[��<A�x���O�%�Z :^��p���
�>����be����?���S���5��*?rWJ��kS�/�!��^�79��Ir�਻� �A�T{�\�fo�g����W{B�#�!#'3E��w<��s��W߶56Ru��-�X�f�|�!��������MWm����Ȩ�6��,M�2ț�I��fr�x��S�<s��]f�\�Ƞ�^.<�Ƹ�$�����aV[���<Z�e�']�x#@?nϭ��!��2�ҎFV��B��)�@�����`�? ��������pWG�iJ��o���\㦸~�+i*�i7dv6p��e�Y��Z){�4G�kJ���I��Z�b���"�8�{����	�9S����(�u�T����d�ni��������ۻ��R�H�����ZF�价Df}%&f@�x3��,����.��Vn�*�5�*���Jo��~!�4⺿keS��z�	V�:�.�\��e�vE��L1V�E;�C�7����a�u�3v��
�߶1#���i��;k��֣�X�� #M㦫��<�ʃ� �6��p:��A�����&�4���3���K�܂E����V&#i��%�H�ٕ�7.~7[f 2�d��.��c�2��#+��7�'�@P�"�NRtu��`��c8�C�ѱ����m�3_s%�Xя^�涴��<s��R2�S��i;�3Dތ>�?`\&�,��Z�`���4=���/�s�nU���w�:G�\"$a�� D���n��1&�J9�[�z�j�6�rc�?���\e���!�9�/к��`�k:hKE�c3��2�R�+�G!�8ɦ�g�j���6�te��KD4T���gE�s��1�//r��|=��W-�"p46ˌn%ؗ�p ����>J��Z�w��X���	�"���4k��MW��d0�x��*�C,u��:[Yxx֠�����^�,�G����~˯�U
�\������	�+�.Q����* �-j�C����Dg�6�VMPρ�2#����G9��� 74�E��g`�H�x��Dv)��+�z��w��ڨ�'o<S<�BdnY������q��ҽ���2}�q�%Z�m����P�ԗ����� �V4k,�L@���'>O,W���#�x�VH}$`�b�[��%��.%3�ERh����"�e}
�N�c�X�̊��~�6�B&aY��ҜX���C8�fIH���mo�&b�5y����$�`sILIk%bc�ɘ+K_���3������S�R1a�̙i��k<#��N�8�I�.�$����$�n�i��K�~���RXA�ݢ�^�H�%�5�Op�������n��l!�c.�3��
�#k�JLGɕ�平��;k7Rj-a�c+�1�G���Ã�b	�K�'}��B1�5ȴ���MiL�����pm��ׯ[[��0��b�*�7Q�k�S!�ȊI��`>���$���tO&��D>W%0�{�Ь�]�r��e4���&�_u�����N����L�$��IB=ViF\Ss4�^���bf5�W⏾�pX�v�T+��,O��9sr*�dhh��vW�D��A槾�t#D�K�K��h���KUL^|cJ�]��Զ���Y&f��������\�����D�R��L��>�f���I���5¦SK�*_���"1��~N�x��͘�|���0�����]�h%�4�"�Xc��>����ѿ�!^3�X�yx!�feS��Ɯ��?��y��ȁ��d5Ù��x��9����F����t�m���O�2\�b�@G�]���G����qo��s�*��w��S�1=+�k�HHm�MN(����st����3A�<(r�I�� �d�Z�L�LC�J �e�wP�t��i�G���S�1�����x@���a'j@Vܭ���L�$�J����Ç�6��`��}"xu�*�ȑ�PF�s�n� !(�`�p�r����7����aA�-�i��@��v+���E�f����i�b�8C�,�5e�q��AfT�IR%q9L�"*��{���P.ñ�V�C""�?W{Ƥj�Ɗ,d�7h?Y%��e&[Q�l_�c#ym��R،;��l6o������ՠ�o�Y�M�����.�6�.�Yԁ<��Ω4kycۓu�/vsVcna9�`��򋦢'���_��֮�D{h�"�ܟK�(�-�7�I���焂��aQb볱]��*�X� ����(�+��F���sE=ł���Ti1T�^xT�nhG�Fbc���	�����$"��a��h����#��S�-t�t�PC?^�[��qe��Af~ֱ�蚸n�V���/o��b�ѹ�^K��h�ʗ��l�0ա��|~�ٳo��^�ۛ�Ĺ�/L����Us�E�0>�Q9g���a�n)���x�Tc�_��(��D�ѯ?��QD=��w5����Cj����Q#�q�� �#I.�I3S�µM��J�� �uG�'�	�7�9�N��ӖW��²U zbo�h��7=N��v�$��犉�[�WǞ��I��!V�$H�z�
@�M	�N��,(Wr]ͬ�U��ս?������O��ɂ���gkD�-iT�6���L���-�L �Ma��8Ò���W��,�q��
�Y�<�!�+�.�C�9�E�/%t�=�7�J���:=M��J豕���ӛ�@_�4{���u�6�B�� M�T��kk���z�%e��L�?�C�aDO���Lϴ��C�>b�%�$��F�L*���1��{�jR�	�pHr����;~�]x?r_�7�:X{~n�����}�lw�%)�����?�m{,�=�b���4$I���@�c�zBR�\�=!����a�p{$n�dAW���8Ha�<H�R����a@k��U�$�����[_��W���<m�}�獮��:8����?ؼ��4��K���^��9:��d~�)8��9k�Ry�ƞos�")�Ѳ�x�%9ձ�S��#��B�6�)H۰�=�!�،�Q��:ߋ�#دكT&�6�~���]����p�0�!�l�-w�Wjt���6���U�]�O�,��Xh}���DgD�Eb�����.�x����.d2K�=�5�~�
����:+O�2m�	�~��o����P�C�Y^��o�(���'�t��|U+���׿z]v=go1��S99Ut�XJ ����)b���I��J�Pz��C3(=`��i%���^�(5Ўc|Q�:L�x~YE�>nq�C2�aV���U���N	���\���<�y0e�g\���e�|���t�����|C�9Y��^+X��
^�y��l=`}��w���!�`�Qo���
�b��|��z�ݠ�f���#(Fl�6qAK��N�c.�)��4��e�-+����Y�/gL �\�Jʨ���s��'ۣ��ku4b����Aq���h�Ӥj
?�ˠh~0���u�{gK�&�X7Tג�����k3��`���FK��7�y{)v]SsƮ���?���z��~����8�/l�h̨o� �K��K�*4z�b�.Eo�y�U=q]wX�a�%fu5�W�v��fsk��w��wjn����hI)���T��X	�1�|�s�� �Ua����|�5�/�O1RN��u�`1�$��ގwr��˝G�dV^������q0�?/yV��Y	@9���2�-d��Kc-[k,� a��:�|2��٫ě�"t�+J��!���d���d�f�\=]�"���;�D������0�#˗J�`�B��u� ���'���<>?S5mJ���>0���#%*.UH�q)?���6�K��z�ҵF0�RT�\;9N���m�G�=q׍� [�v� ����Hٽ��#�\7�a����k�.�����1����>�u�(�̋�0�t��g�XH�D^%�Mɘ}���1 ��v�ȮHz8��.E�:��NU�=#/���Ơ�JC&��k>�-�z���띱!��?~�-�H����a�3fW�Ož9Ce��:`��[�}g�I~�"��$���jU��r�&��Ͷ����K�u��K1��>���F��K�� �3-��_Up��?��d�qD��ޏK<�gf�a0��h�>-�u"�9�[R^fv�X�|�F��հ�'Sh�����K�k����e���&v-ʊ�8@�#�E(U��}�۞?2�+I�5tA��C	Q�R���Yt5\�)��d.���Q���(�6﯁�b$A̠q �!3�聛p���O�fVT��9�u�y��n���aRS����-�<��4��VlO�"�e� I��7X��\����t�&܍���uy�A��� [�	�˛Cp�W��;%f���z+��7�}��{n��E��D�`�еj�u4*ɛ��"��+<7$#��6��[�ʥ(�bg���"ik��v��m���>���4����N-qĬ$Y�������O2�+�!����t��!�FD�Č7y�M����m_�l�ϔ��s!���y�?r���a�08"�����׳���h�%�V�	�"����.dԽ3ZZ�Q�
P����Ȉ����Oe��IklP�Z��P�2�?ٍ�M�����lL�yb������FK%i��� ����Y��u/�O���u��ysmT�͔wr���ڽ��reĪ9�*U�&��j�:��óF��{��+S������V�<��Xrp�X&E4�36��*WRSi��:��orJ|�6K���2a.df���g��}�ź�R��5�����PiX( ��4#v�7h�=��1I�MC �U��7�!�NIB+'�g�J釿�>Fh*�P�A�(8�9.л݀H�1s��8)od��ـ�����k�O�*�w��QZX�x6�E��@QZ����>H^R� [�z��C��<�0�c���ET��X��=X c@�m��D:Ѿ�������yl���[^!�@���Ö�4COR�J��f���>-�ɯ��'�s�����@�C��d�����)wXa��i4V�{��ӷ��{�o�	9m[b�@$H���q�r<�C݁��FTW��l�,�3}?})� Ew�G�-�K{��4ƭxc���Tn%���qE��I�D�"kO�y�q��&�խ\����k+;�lS�J�2z�k$�Xw#Я;kORUvab��H��J��ao��{��=[�*U)
�i��g����=s�q��px��5_�W�G��b�=f�)J�3['�O�"��&�m?WZ=y������L�E���_�0��SD���h�`��E6����H���c��]�
C��>Q+_��T��@@���p�������� ;ͭ��6�xt�;l���Ui�}/�b��NF�|��8�/���mf�o����w��ӽsw,c�[����ݸVk[Lۀ�>�<���7�HihZު���&���#�2i?��j2b�^@ޝ#t} ��`̈����/M/)�~��6�k�ⅶF�ɍz���?����$�4��u�~�ɰ�Fhe1	&^���N;�30�%-��e8?�K�TgR���B���m��89�c��N{�y�轐l��Q���y�f<i��L�ה&#|��`�ET�eQ�v�^�#�&���<��Jf:�p��zQ�BI���'��n�Ƿ'Z.�W��<w@�"Pv~��Y!�Ѣi�'UЧ��R������QG9����o3�]e&#:ó�.�o�O��������\v�!��5�8ZS.�{j�'�P��h����%2{��B91����\�k�M��>�{�����e!�p 8�����2�"/������f6�[��ݙ���)�!��.7.|j��͔f���=�/�!Kͥ�cD�g��
�@�(,�E\C�h���M,��8������M�Ld���'ܙ���& �#nzHTA�m'���Oxi��s�M�m�o_�@�@-�K@�I8*ir/6�굯:d���r�/��ceI
��*3;� �� F���%�I/�=1Z'�i��CAjX#�����];O��;6o��&T�0���;*�q�^�20r˄�z��d��gF�InZ���bXbG<�q��"r�A�f���b�5R(a��;Ȝ�%�23��OQ�)�{/���n���Y%�`�BK���G��P$��, I�6+�縼{-DZ�ʷMɌ�I�B�*>�4�#) �z�M�v�� I��%ھ�Q�|��rA�FK����v2���'I��z"6m��k�%̸�J��V�F��"���^����W�t��P��BE����#A���cp&���$�h�[?���׿�~�(�fv�>��l�{M̴۠(�FN�kPw�&Q��5&OPA���?-�[���u+C����o�n��4&��w���h�+&�:1WX��냥`E=��C�N-���>��n�8��q���{�6A!��S�D�h����˴bd�&��/g��ǻ���'�gJ<���xil�c�Y!�S�S�#�M	��8<ek �)��H�$��L�U"�R�^��ۊr=`O=�[�2�q��Q�	i����F���#�Lܔry~If��cq��e���fT��@�F[cj?��q�#cE��x���]4c��U�Mu��s�g��|l����b��;�l���6�����Av��4[u�V��~R9CkY���8�`G#�g�"dw� ����uE�z��=�9k.$ـ���d�t:X8�8Tx�S����g&A����g�1�T���X�	���A#�K�Ҝay�-e��p�?ċ�
!��4��/�� p���4��UY�JR��R&��e5T�e%9R��]������vc�v��I�i�ل��Hr��(�҈>iy+���	e/Xh���otE��c I�u6�"�<EX���够F�_E�a&Tv9.��s	9����v�ȼ����RO9���ɕ�dVC������+��B{�YI�X��C�q/��=�f�2�$�^U����M��t��1Z�`Dx#�)������
�9���9�������F��M��!~r2����j��h�n����y9 ��I��F<� e+ʾ|j��wo�:5+�n�.��1cT�U@��|rdl"�/(����xF���\�����l)	:q�a��:A��\j4�8��畲[�X	�8���j�~�OkG��P�Qj2���K�/��-&��˔�
��d&�Z��+��z����+��ӫ4*u��pɚ.1�W�3�i=�Q�ao1`C�	Q=/?Ԯ���7 ;�:���lK��Q�J�9����R	 �_Fg�9��ӂ��Tcy��W2]�d?c�(*
���y����ru�fԐ_at?��9+ ��%)���9�(�/Ci�C5��	I;h�����C؇:���fgt��=[+��#��}��,Z a�v�]�KLU/}��.��,Я�`3rH�
��e���Y짉0�V����hOQ�)����NE�bw��M	� >�Kc�u�m��Ě�
%Wo;��O��Z�\G�7l�?��g~^&�8�E����K���@��#h�o�5h�d�����O	���b�Ҩ�0�t���#�A���1%9-�����x~�������R��_��]]$��K���vcj��9n����G�_��M�g2��җ�|���6�oh˛ɫ�M�|-��ix(2�[�:�N.56�^:�T����r��?���Zߚ9�m�{��b�(8ۮ%F�q����>���BVr'lG��z)�����	*��Y.u�b�K,�诊�����qЍ�M_��֗)�f�^�g��eN�ذ�M:D��{v�vW2o�Z�*>Mn"��/���@݃�z��N�>��괫(o������4L�4���r	���^�,z��J��{A�{� Ruۂ����z��&��ܙG��*�@v�mP�,��B���sH�EJ���~�rS8��@��cr��J�����ͽ�(���&�y͓���:��͡���y�[���
U�۰�b>�tB��	H����`��Y�fъ�r���^qIb��v��$/'�C� I�C���D׎�lk>_9�ۮr*9_F4��R���0�+iyf�اP\Ĵ���FP�=vy�F�Լl G}Y��X;�5�G@B��
 (�+<,I�Z��k��ǔD]��E��z2.���[0�Ky��ޖމ^y~ ��!�׷y��0d���=��+�d��L�)j͘
��%/��w��^��z[L�nx�C��'x���s�!lg:g��¢َ��� K{M4�\u�[Aw������v��re� ����W����a�<��B��,`�I�Po>e^/g�9Җi��C�I9W�^ب���a�κ����������+u�p��� �/������Wu��E�#=�c����+�:a��s#��;��)6~�'�<)A7�q��5E񊃕��֑<�mG�čF����m�j`l��� ��5Ɩ��$�G�qt�}��!ZU8��̵�%GŪ�%,���'�!�)ң&`s;�'.��� �pM�'�e4� �5�gl�M�=�ߌ(��Eس�@���\��K�p[�����u�o�aF�́.�π�ԤP4Oo'\y6��I6�~�>W�1q�n�/�-�yi�{��}nE�ۭT��V/V�R��r)Z�Rf�x֯v�,��V51�ᶖ�"/�Y���}T��{VCaA'u�
%ьY��#��n$�s��l!�+�W��	(i����M?I�7�g<�\	k��Y�1![V<���&~+����ǵ݁�;b%��}0�%!=���ܳ^�� aŋ ^- �.��L��c,�x~�1�_	.��t[��4�(�P��;y6�B�Q ȉ�9��;N�v�h�(s;�/�4SY�����z1���`�-o@�������Km0s�q�*�6�qg�Yڭ�KE~kӜ�]\@�۶0���IL�e�,����_�j���ɨ�BJ��H�'�+�l^��	��ۖiT��f�Ώ�����lY38l�b�o϶j,05K���]H�>cR��c�$�t�N*��؀N����B��Qԧ�螢ڼA����T)V;	oQ��
�8�Yr���w�x[��$�6'7����
���xZ�Sg �3����GMy�(��|�7l��
�s��?|l�xVtV@;r�Y��̨Z�$���N����U����(�exݬl�.Z��p�Ą-P�!W^`��Q�E���;
�Б�b\5z����r?հ�l��J���5�7�m0$!i���_��ߠb�]�\����#�4�$"g@�5b��#�Y*H���Ϥi#�;�|E_t�jD��zMؙ{��� ;���0L8���*ڠt{��{a�l���>1�"t��2l@��[®,[���'=r�*r��S�B׫$"Y8������4���τ�I|YS��]�� �[��54��ë��sV�PG�Ũ�Lj�:���w'M�Ӱg��3B�[#���:��?�kN������)M�=3�Đ�)~r�U�iy���L%�~-�8 =Z������������s��i$~�
�����:�@�\���**z�����gC,鱋�������c�*�*���r�i�ne��b��#�z��A�oX���,�~��O��]��m,�{bs�^8�<���O���W�B7T[��������m����o������q��H������ksS=�nt�@8/ �8���M��Tc�2� �(���gk��	�411ݻ�r��]4�R3+)�V"��m�T.a��I@�"�����xOP.r2�+��=Sk�"D�$L�~��ݟ��³+
;�)�)��k�mU?���Co�2��Kr�oB'e�.R୩�Y�?�W(z�/�dj��U��ܱ��-Y�������,>ڻ�g�Uq�/��B��̒ߩ�[$����~ĚG��}��q��J��S��Ю$�����]����}�f4�M���͆``5v��4L~co�J~1�I�����a��<��evD�wV(u���x�΍U����������`	K	=����>��y"�P�3Q��7-�ĥ�DNA�A:5Q��2�L<s�rܝ��WptOZ�3�㺽���+��2C�Ez�K����4��_�ӷ��X.@@԰���;�o��
�"���&9�H�2.�=+2�q�f6Ұ����b�{�(��V�(�&z���А�ct}Y����e�Z������`�@�(~���LL]b3t#�M-:i@X�V!nx�e�����*{�D��-rAkp�b���3�S��/�������V��HG��z	:WsMH�������. ��B�͊��8�|Me�v���x���æ�C�������/l0}:��]��N{D6,[��n�	0'g5��Fك+8lL��&�-�O9�ɬ�i�# �pl�[�u���P*��x��h��;dM/�J�4"��A��־�{��_���'Wt�=Lm-5拖�>9��5Ԭ��Q�w�v��"P�øQ.������ҵ����9d���cw'�P�r";J2��Z&�u��.6-=˄XP�Q2����WV5HK��B#����=�-��}Z�,�"��<`a�*�� ��������;��6�~q�$maK���3�b��Q��D���T�hރG�'�|?k����*�T}�G,:�iUӨ��c����:��=�5t���I0��V����ky#�\ah���pp���jH����/��8 _nTp��S���|���箑^[����4-M��˘�&��۞�b��%F�Q��#�I?O!<|q~�{p�ʗ_W]�D�3Bي�)�B9���K>�G�i�<��햏�����i�x�|�X��"4K0^:R�|��u�)R����/hv	$UHIPًh���^��-0}5B:���|�kK��nUL8 ��1�Ʈ���6W��[V�d��2�_��W��l�H.��B����� Jy�R3%����pQ����r�V�IKiv�U�;�*UMkޡ���{6z!e$ZF��0=�ȵ�xܣr
v߯����K��/L�vEF�J�����M�Dv��}��i�G�v?ׂ���ߏ9�Ӗj2���nNv�K$>!�e�0�^k�7��5��1xCƜ�W�YӃ�(�N9�� k�fÒOA�h���FI��jh8�� l!8q���e��ڹ �@{����^��+�MD�g�`�@;&�0��)�M���z<u�bɻ#Qwk���Ꚕ�fQ�p!�'!�����Lá#�&�)T�Dre��x��{"^��Z�@���ǖCzp�����c�C���t��q熔�s�>�#�C��O0�<�>��mL���P����l�z���B��d�J�
zvX���9�6��]�
Nڻ�xc֕����?)�,�j�C�+�î� �RA'�-.4F�5��"��-�j���r�r>,<�Nk�1�%���O�Z�w�k�`�Ȱ1����\3����!��?3�B��?��R*)��g�S_��4U�`��pz(Q��}ꨂ_�6G2�%!**�� N"	�W��)޽��^bY���O�M�dK� �R͌W����2��Ȗ�$�
��3P��d͹b��ڗ��
�!wݦ����@�vw��NH{yV�{#p��(mTI�����^-�9���`��[4�Q%qd
�®�
���Wnmn,��3�(X��uBGh�&vt.Kn$��0��j`4��#�������W�Y���U(���2�Z�޶!{���y��N���U�:�e���3���U{N�	��m�--�is��&\i�����m� ��J#�\]��@��=���mb�+Ձ�����Mf�ױO&�T�y`�W��]�)!����v[s��a8���U^���r%��e�Y��&�[����y��4�̜�!����:��1�T�Ḿv��~0c�TR�?���Z��s��/��z@��BN�SK�	�ޑ���G�E?�����ȝ�IB>�[{X:�|�y��B�o+^�#�0��M�;s�jf�z�#�->�r#[2{e���i��)�t�ƸM|>�$`H����	�~Y܊*��M=!�ȉ?��'�@l�w��$�ٍ�	8t����UDК���ˠ�*9��1]�$K׷�&$^��'4��4Յ
O��TC˜�P���g�0�;�y����K�f��`�uo��)�HJiXNw��n�B�����8�6�5��n���k�R��|�d,x�w�~�]��2��H�z����t��WV�#��8��D2_W����M�k
[j�я������1�'5n!?v��&�������c�k���zk<l��7�4#�p��`��3���]��u�{�9��T��p�G|�&�>��c��xGi�	�	Ơ�ۢ�\NIB��<������@ۻ��9�̿e�5���9��-i�a9U��Qȇ�W��e5~���c;�-}�OM����3�
�u�U�R�V��*yn��Y��>)!\
fK}��O?�2��G�����d�e�Q��IFQ�ns��W4�ϳ�@�?KVAf�5�9[홋�nU�oȴ�g��*+�Ij�϶�3n`N�dĸզ���K��~�>2Or9L�ao�~�`8�;0`�`�m	=�NeXv"�[B�
˭2u��JZ��#%sn�NƏ��/�hz�p��X=��7l��Hq����'5k�8쟫0��}%��'{mp(7[�6�+�<�6�?��8-����&s�}�w�������{�S��@�J���+�x���@u��D�߾Y�$��%�?}5��xA��pkg��eB�_9q��y���
���h���د�es��Ee�ͥ��>AƆ�;��Ҝ#dk�9 UӋ|�� ^�եƿ�%*�C+t�Vai�}�?��j!꭭� T�~�)	�
�1Q��c����r
����?р]dN�/��q���X�5�cMm�H5��z�%�o���[�nq9��Rc�y�l�7���e?�BN%�zz�y���W'<�e� �=g�A�p[)%)�+����sW��4LH�`�k���6�=�j�����*���2H��	nOIl�Q�߃4j�o뼛"��G�:�K���.,�g%���I�n��ú��YN�3�>4τM՛�U��b�A���(����;i`��	�dn	*�]ED�@@g�o�B"��"_+UG���2e2�8�"Q:�&�(�T~�����ԓ����ػXKJQ*E�/z�%�Bf�~��r1@t'�\V���3��H]�a�,��b2��t$Vv-Î7���^���h�W�������kpܣ$8�L�EĽ*�d���.�
���c`��eXi�����CΰD�}<gm b��t�0\͡�#2\�.�����1%a�& j(n.X
�($���Tm8%�ls����3�b�h ͧ���Vq�McaZ<�����L}�E45��b��zzֵ����3꘡��s`6�`�ϓ=�\����ꛉ��$�	in@��m�.��
ה�@f;c=�cN�Ӱ�T~%7cKo�#$w�T�u[��ѭ~�ct��$�0���a�V�3oљ{H�C����wK�G�|yY��@v�����k=@y`����D垭��/ J%|[�8�{�:~�Й���M�M:�k>~���mѡ���m	���$Q&�wr>P����ý����1ܬ.
��Z��-�fs%\"�d$t%�]�Tϵ��}̓�by��LIV��+�;O�-͡!��֐�*�z��S"	?q"��G������)�Y&�n��M>/8��+OJ�c�"��^+@�j6EM'��(a=�񾆻�溾KmN� 7����x�KO�D�d����Gp��s�lF�E�~/�	����,�)����\|�pJ���}D�(/ە�2��?�l5����@t�!���_�vk-�S�!g¦x^;�����,΍K����ʦL�=A��jCHR}� ɶD��(wŪ�b�D��֏�:{h&���v �VLƖ��,h/.�U��F&\Y`�~HuM�$*,)s�f�Hk\�$w`��Ѐыo���%���]����_��� �R�V1�q�
��|�TA��O	��t%˄����9JK��)a~��(-������q��ȷ�A�gn�7>���2�%^�5|����)��m�pÒ�$�?Л�`o&�ڶ�8c� �p������#7ƍ���+*鹝�[\�4LC�����C&4~��}��I%�����z�J-̽;%��W��v޶��d��t��U&말�j-�X��{�+Rq_�$�@���� ��+-M�+���&� �/��E̎�p�Ǩqz��ɓ}���m����|}�<&�c����-@���*�K ��8 �*{?9]��a�M�Ӝݸ����7��l��Phj�R�BF�$��v���n�����!�
������*��W�;��#������;�ҕ3vB�)��4x���m�o��y�N���2  �?� B�]��m�d�*8��6�R!�?siL��*y(x����t/������=f܊:O���ٱ6!)mt��Y��f���M?���F�O��V,��(�|��Ri���F�;�����e��cx X�W@��aSS���=��#�dd�ә��@@>J�,���Mx2˰b'n|x�[�q�7�鐹@mnG���2�b�!�$�@ne���@��L��	�"A}��J�rӺ��`Ҩ����17˖H ��x�k{qEo�c���-H��J�c�p�X��d�=�Scp��ğ��������B1�_��>>���Jx�Ĺ��_ �����M?�r�fj2˫}ڿ�H���OaX=O%��ۻ����M�ȧ6�O��i�|�� V��ԋ��U�����"fG��SKMz� i�1��,ԫ��1}��f��������
�,Xk�!��@�E���m�J��`j�Ã�H�o R�&�ڜ�@�\*�W��J$#?�	�|�:n��оg���{�K��X���=����H�R.��*�����ȫ�:���9�9���xIW�a��o��U��v���-�n��HC���;��z�2�[PU�9(���B@��}��)�Ye]���@��f(~���~1�9�8*��_��8\-(VM#����Yn�(�b5N9������MDPb����=�8��D�/��F3�"�UD����HGX>�@�����V�$PE_�~�5W����g�IT��N��C��P'�U,,^ ��u���o��wÒ���E�a~(�e3�<��Q7�xQ,�~�����Kyד���ڀ�
�>�]��DXC4Q�������]����_C�b��'b�N���o�ӪZ(���M��� 
�)c�	C	 5�<��p���r��R����A�ENh͡*��N1��Gxy+����L΃֓To�ʻ�|��i�h�!��y��ufmT���.�C{O�Cĉ����ea o\�I��S�Ԥp68/r�D�bt��u����g���|g���w��fK{Ҧύ�i����"**��uǧ�4�ኪ��D��������	�X
��8U���hŔ%�5�%�,�z���J�A�'9�pe�g��KoUx���8���>��_(�Lcx���1
�����JSK�yǊ� ����յ��,cu��H�����E>7�%�8��$]~n�ZsJ�%�"�(�qꃲ���$0�N������}@L�@�#�S�����<�y��*��?�Ϫ�S�U\J�@��J{ê1���B��1�,ĭ[�ͦ�5�!��V�X0���6��2���������H5\�=I� o�B*iD%A�2z}X�|׽L2y�	�[�1l�N���"C�(��g{����lGZ�nR��Ӡr�rr�7p�B�z���}�A���ʉ��+�����\R��"S"F�������A�Ru/H��矅ˑlŅ���`�����cw�E0ްK/��!䇈� k	���GMƄ�򓒰rq��_Wa^p�7󖂩��49\�&����:O�/����
�ֻ�����Zg���}״�{(8���:�5�f3��~xH:��������ʱLl�o�"y[���3O�s��И仔�Ahnp�n2.aH	ط@�Hj�F�������7Ѵ�
D�n��0{�\��*��c���;��7��P�u�\��3/�{4���D���^��ˈ�a������ǭi�"tk�KKP���z�V"a4�m��f]�a1\�����*>3`���t�}�͠o�0L'J4��Dk��ヷ f�9N���+	3̥H�谇�q�8塁�$��[?9�!Y �XCm]N��h�����i۬�ޮ���ҹ����I�Ǝ�gg���k��.�Z��x�ғ�$��AZ �(�Ȩ�ż��4��2l�3K��nI4�/�s�ș��͝�R=�^��w�L֕�47��6�d���J��q�W�4�ӵF��A]�T>�	����!-��^'V�z��0��������h�睈UqwC��I�LU�Y?�J���˖�ٍ�J:5�ܻa����۲�G���k�\���:��Պ���J��d�l��o	��
�nY����(�l�53�5G�A��1�>k��j	��f�����ny�@�\~�ِ�G`�N��<��[f�٣��v�$Z4D��	x��h��j�p�d�Lq�Sy~��2��&���nd疡�U�
����t�(D�H�+�D-uˣ��E��*�|ϻ�l*���i���:����PV&<B��p|�<�Q��֍��\���~.ŷ��/��g�L��!&��kR�q}�ᣭC��S	P�$�n��t�#2�c��Bi��ͷ�J��v�9wq�Yd�0I�`}[�M��A���jO�r@�(����6�H _{���0�#��i������>%�3����.������.v��"	}z?�z�~�<)*R����>a����m�%��xSSB9x��F.��%�	S'7t��z2��ޅ��Y�w
�`П5m.�mx��;E����Qn�_�>w��mI������i�2]k�G
�Ιp!9]��ZkA�:��n�epMOŵ�4Y�`���ʪsJ�����V�Qڛ#Q,.�cm�x3s�P����m�P��!H ί���ɱ�fi�|f��e�*#�S,���;�k��5:�^�	�T�STHY�v.s��a��n�'`A1���9�
���viL]�?��S-9�6����zV"o������G��ʸ	�E!��k��>Q9.j�����(���$���s/*�Ę4 ,�Az���z�@��#��O�S��<�`���əDk�T U��Tl�7���D��^�６%b{O�Z7kf�x�
��[NC�Zclǁ���8��3�������uQ	 �x
��B�����T���J�����!�RM�e����j	>Ă���%U��0�[|`��������OzcZL����.0Fc���c;0�2������ɍrR�Br�Q�ؘ���-y�8�<� �"���Xu�ᓑ u���G�˜)��E�{	�gW�m��j�E�)Pw!e���k��U�w'����='hjH��+u�&�x�M|t#�k-�xj� �Ț0@��3�:mE�E��/R��B�_.��@�)�?7�������d�ز|Po� ���I�M��*'�TZ����U(g����2h��c�?�V�џr�5�V֜V�}۬�F��j�z�ʖ똑p;���o����4�/�ʾu˃G(P�Z��X{�;9�͡Ģ��w�F� sUJ鋾*�)�o��hx�[�B�vA�����^�7aj���@�4x���` �y PYk��dRMZZ���T����:qT��J@�[x�X���$�Fwv��*�>�c�6yhr�㢲�ж9�e]˺���MǬPo^�'S��D.7Z]�p��Y-t_/�msB�ɳ�_y�3�h��� 	0Z;k� w@((��C��$<h2˜���=�d
�F��0�>l'�#��풋��I~�Y{�����/=�ApAj{:��&�~7+�����6��񣾶'�����7��	��2n�bW�7wӐ�E?&�A���h���Ur��G]�f(Bŧ%R�]�@r��K�9�Yu~�������v�/<~򍫳d_�H��L%y�2��`�ZT/��q�g����&v�[�z��2�^6��`���&��A��͇:D������z��/�4o��Ĭ5o����4&�	��Ҳ�f%r�-}z��<|��O{檥�e_��6>��?�����ԇ$S�d6*��
ԭ�^v��h�0
u1n��������7vPO��<�C��Lcq7�@��U�������_ 6ֲ+�K�� ��\��Ht\�<\��{4���a	7Թ��Y%[���oWhʢ7�A�'��ƄD|����^yWj��z��M��ױ�4^ℙQݸl<4O���. :4�]Fb(P!��RQ,F����>��|�k�i�m��^UqG�@�e��m��'�o[���>Y�ߙ�I�Ǹ�U��BVB�ECf��8�\�IW⣂������\��S��$*��َ��a-����O5�#��t���>۳A����V��i�	<v�:8v�O�J���y)](G���J�Ȥ;��d�}��Ϸ��re����GQ��%
�c���	e�O�� ]c���v�6^�VK���o���(2DL����
����K�����m��}�D2L��1���xyp�'���n��}x��[z���f�Mep�Jܠ��MD��	�Hk�-�T%��k�����[2�h����C�c"JY�˶�d���������n���V�/�`��mf�ٻ����ȑ�X�s5�%�d5nƦ;x�U��<Wg�/_�-E�r�1��9�e�`Gѕp��\V$�cP�\��}��␜��{��p�{eʎ�v�DK�����(�,�r��:#��P`�Avl��wu����J�8�w�B��i_�7�e&��Zꏂ��}@�����/.�WΤ���d��5ڦޫ3y�!��a����S��	t�'��Ye�q�F� ���w3ف��	Ky�n��a���)���$���eL7��=�}��D:���i!E;�6�{�G��|��ϡ�u�t�I�˦���&�FM4:SӢ-|�J�c�0;��:y�~�h6b��RL��<$L��H,�� (���e����&hb1�x��6�S��ެ�L#\,=3Ԩ��\n0���ܶUēl��	!�U)���]l<>��yw,��H�x�褫A��;c3�����R|IG�mH$�V��"��xu�9�^�ՆY+��h2�]8��ģ7����]�;h����.�B#�%��We��`<���]~mV��5^k���B5�_=��s6�����/}¡7 BG�f_��у�3���а7�=L�l�fצ|�a�����O-�����ƭVn��n�L��"�잕�O�'�*�2�^��h�3'#�qm�*l��g�B�E,��s��]�)��Wm�ѓ�:��\*Q?��A�V�~��+��~�K{):L����:Lȳ�sWS��,hǑ|kRT畓ۧ5��l�_�gܝ� =M6�
O�1,H?���=u�?HӖ
��^N'v?-f)��[*��&�,�Gb�d��⟺W
Xߘ���>�.�����"���B�	�cN��o��r -��u��]�si�J�Z��D�Ō/�)2�~�a���Ї�5�b������å�)�&vQױ. ?
�pJܖ�u�c�홄�S�յύ��>\&u��|84��^f��\@���MŮl|^5Y�}.��+x���y¢��c���=!��0�\���t��ӟ���s��@�/C�6�y�>��$����z��C�t���\/U����$#j��+��x��˷��吔i�9
�s?���|pNi�����I�Sw�"���Ń�	��N�y<��o���͠��.�@������oS��UU�	8����t�I��f�X-����A5`�� z
�3)H��[�,�/ř��}��� ��"�ʄ()u<}�����A�-�K#����i����"��0��g]G?�"�	b�!��d��t(J�#^K�	��R���{@Q�!�#"1�����-i�A��c��Y����o��9�-������S��yrv<x�ky� ���7X�i��Qx <��u�N��U�]us�� ����I�)�ݏ.Z6j�Et�p�vD��&԰ĽzN��7e"^�\�n�f��@�5��:��-����ذ�w	D�f�+Iq�l�Xx��(���_��3��pW���TY�*��Y��[���YO4�������`��Oq�Oʞ03*��@���j�sb��\	���6Lmһ���YhZϼ�.W��;]B�����
X'��{fB���처��Ƞde�~��b�jL���s�ZQ�E��x-��|��к�~����.�|Gn�7��g�a�����7�2R^��А}g�e�qN��Br�3�ɧ��څb6F1���KѾl�H�Y-�N:x1��LqU�I����oSZL��E� ��F
�93$�����Whqt�	�| ���gW�V5���;-��)C<��h�����s1<��#�Է�ɩ�ek�	��'�S�7���!�m��ިb�;�	F�ž_����D3���	w{j�% ��2YN�v�??pD�}������4)q�@���M�<Q��.�� �����J<c&�2�o�܅��U��wU���
���u$���o���+Ne�Ͽ��!��k �~�ϼ���[B�s�l���8*�S��J���kn��5�Zũ���ǖq��� ?�哯��Eּ>#��+�%K��'�8J2����,�`|���E�$�ԅ�Yz��
$q9�[��$e�k��CN/G�T�U���Rs�p�F�[a"�-ja��c	���q�J�E��e3��n�g�y7ٺ:7%�s5�˸+�ʘ~0��W�E]��^� ��V1��)����x��"[z���kt��F���*J-�Z��m��F	�ia�O����B��T�Dn�����%̽~٤+x��mt�tU�]e�SF�!���r���2Q%�q���K�9'�	Cl��iE���0[�z�3���#�5�60��.�8!\�4L,K	W#���H�,��t�����ٲ��x]VC�?�A�
��R�u��	Yv������So8��.��L!V?>$ܹ4��){i�KH��\R�b��	:�#�U,���zv�<�Z��:яg��clg��?ކ�͓��2��2]����E*%��I�8��Kd��F4���=̤�N���Hj1Y��Q��ފ���p�1;�D\�h^IPvja'X�Z��M�؍>g�~���?�7�J������Z1m�}���E�T��hu�/ _�5���d�h�'LP��+��Cc���K4ky�$��Q �H�P2'(�u4J;����q�
b�������)M��ȢLn��x���xʄm�H;z���s��
�΅�U�2�&��p��n�Q��e_Y��q}E�'=���s���[���UM�F[���A�Lc@�`�deݽ���(��Q�7��)�UT��ƾ^�Z��iwW�1y�T4@�����K��.F�����s,&LL����k#����?N,��Kx&��C�b����:U����=�TXa���
'4���q+�{%(�D*�[,>w�}�f�<P� �9�9Β��w|����cw"��Ղ�xf�{ս��L;l�e_M'�W�ӻ�v%.�u���+��P�9�~�Ѵ���<ozk<����b���BL�b+�ΨB�`��� !2~�K�I-�డa�ɱR,����G�����2}�"�\�;���N��!�ߵ�z��؂毟�L�O$P�;'�(	�~����3����D�t��}��>5��b�w���j�R�q�3��e�,|�JJ`�=�~�*Ӷ���g�x�I	\FK"�~�<
{��0��Ӵye�K���
V�rT�Έ�e^�F{�9����
?Ӎ�U7?����z�]�f���,3Tք�(a��n��L���x�&���b�����ixD !���#�V��Ӡ��z+:|��4S�%�b�'��@�m��W�wҚ�O� Y�J�WJ���=�%��5]�k -7fz�>�6�H�{ۢY�S�D
]���b�^ح���F�׽���_�ia��4�1%�E�j)���)& �Y<"�f�# )����Go�R)�A^[\đ��Jv`��ַ̃o�▔gwߑ�mc0�T�91c�!i<y�]l`	}��➦p�m�׵��Ù�?�J�9b��NQo��|��kI�~�d~��
P��[<�{���;�s��Z91���ҋXn>��ns_-�_֣&s^���~�
$�O2d���ѫrE�)L�d��$� �K֟8�(�P���@����������``G=2�[oF��	_RL�&��IS�*B�r���%���~��PKl}﭅|��"�G5>zN7��#�û��d4�ƗW�0X��T�y� ����8G���¶�׀�������^�m�G�O�*�Ld�����y�@L�(`6��bj����5�*�[�r�!�{��U�ˡDg	���\�������nҞC��Zk���i�"\��j��04���پ��8�L��}��m�pw#a�>�2��܅
ܘ#��=iz��Af��Y�����ʔHfF僻^��p֙���� �t�%T��J��t�>#F���=������g�j���-���M����(1*�@�_y`2�v7Br�?ڿ��!|j�N�8^�����^��1��
X�w�w��ܢ}����̖�k���)�g9������Rnڍ�?U>����\MF$�<B Au�7_��l��B��!@x��v�U�4�[:� 6��ѢIa���k�#���X�X����/Ep17?W��<*�C�Ayn������x���~�0�c^���X�-�M��|ø]W0���Nz�뽥�ڎs�jq��O�� ��h%�����
����wKK=���]Z'Ւ���i�;�3/����>�0�V����ڢ�����4�>fi�C��ɪ�5,��f��8��D>@zT�p�u?b�:�K+q�c��f��{�����%W��/4Uj�Z�P���bG��%b^��NJ�@�1��}v,m�nvg`�ߝ�e�(y�J���}����(�V�ˬ8)��z�ɡҪ�`�Rݗ�Ɵ7�l�M��?�7�76��p�g�x	���~dҺ�׸[c�S�Ę�`,�m.�HEd�@��m&d[����J������=�н�B!{%x@6�e����&R��~����q��}�[Y�P�q�g�k8ߐx�=@�.�t��uH���)�e-�V�9أ�y ���r�xa6�I���ԑ������wh �-�>i\��m#�*�$0��J��Q����@S�\��W��lČ|jx�%�jD��\8nw��]Iq�0lcj޻ (��t�S(H������赇��rFRB�L�v��	!���$��ٹ	ӀK��|]�l� ��u#���GK��W�q���]!�[TK��G�[�c^��I����j�O@�S:B�J�$�x�S���n:	�m�Su/����H�.���S�d�J��>&��QG�/"��WwGdfCk��ڬ�W�P|	J��o���K�x��5�?#\�x��GF)���V��Hq����|O\��M��El��Nŋ���2� (KLfWj�Q�^+�tWe�?P��V��tÛ�E��+�T��)�"	���^1���`u�S�2�Mt!y?]2��MV�rH���#�n��І*O[N��V�܏�nh�w����s:ťr+�I%}��-}��l����y'9l}���ě%.�vc���G;'^t�xIt�?�d;�W�j�ې��xf:�g;���)K�ߍm�|O2�X
�_�T*�;���[̦<}�V� ����!�A-vl�e�\H��R]��`*�_ß�ɡp���`�6�3`aqݱv�N�N�iV<���C�L��\��|�k�m��m9�TªR�\�Q�t�U��� ø�b��4鿭c��M��=p��7���U`o��RMN���<A������K���?�}2g�ݥ��@��Bl�&�X�c�vw�w�t�I�s�Ç�����Qb�9%�D�a�y�����j�;������(#@�X#G%|ej��|���͙S�o�Cd�����nLuGV����"E��c��}��h ^�e/^E�yX�{�jK, ���$�A(��^��� |<��[�~vi��O-N; =W]���_�8;�Ke����]�ŋ���D���d�t�j`�3�_�y�=�?��b�c��3l&�q�J�L���9A�}A�${�,�oTK*�6�HQjA���,� ���4ف$��vL�3L��ҳ
����xY9�W��l�CُqH��њ�鬾�9Q����/������DHb8	EnR)]Mk��2���inu9[�a �O(�޷8r�;1�R}���B(��3�� Tr/#����lֻɌ�*'�����ַ��E���UZzi&v�2�]\��¸j�p����/�ʴf�,���'�a�b(6�7"��.�7'E����E��B�B?-��_��؜	�n��ã�㳽�����I�0X���@�4Y�n�&6r�6o�l@��X���J��㶰�zz}�x�V�cZ!A/l^"Y�_�a�B<����TK��oq�l��كݡ
s��֘��!s�l OY�m5�.��}ðHwC2��!���vӁ�n�AB��h�[/|�,���4=�w�(D�X|+X@�����H����CA�K\]7;��H��|�ʺ��0n����\:���U#�\���iý�60wK"�|��g,!@𒜿�S���ê�4�.p(52���M����c�B������2}�\���ʅ��|�A��CD�J��X%q^M��Ƀ�^�$���JR#��tH�3��7��ɜ��baP�je��� ���Z��0?( =�ND����6"�8�	?�xἢA��XCqc9ڒ���V�Y2�t7T=�@1��m��_eUt<�À��	������S��BI��B�y�2JJ�H�Կ��ܝ6��'̹�M��Ƃ ��%G�Q';;������r>����'H�$��Q�$�8�7'�|�E0vy6���5�q	�o�%I�d�&K��@u���~r��P�3���\�q3CH5������v�~���O{�o��6ۃ�ı�x��1WU�h���!n�K)_X��P�S�·��%���0T�w�|�|�\���ΰ��H�b� ak ��wS{pɓ=1WMCu��<6��Ճ����|����Vhr��Ƭm^
FjG������7�0J�>`�f�ߵe�ĵ�����r��h!�K���� f`W��l̃Nn�b��
E3�Lb��M c��ߜnZ���?ǡM�y�)誰hG�<=��ά�c	��0\i#l��r
 ������k�y�2��v
�)#3i�9�g0��_��cG��m��}�4����jqA���ҩp;4�a
�j��SQ=Sy����j�T}}��$�'L/	'p
+F�C��qО�F�!�Aw�u�M�}�V��A2H(z�Z�5:^�3�w�hĿ�S��^��n2�~�1��i�vt��s�Jl^��!j���4��H<��}4#�1<��zX�䔴c����ȇ�Vi�I�%�_�4'�TR���V�n}���1��s�W�/)	K .�o��pxs�*�,+�H;��b����:�bn��\����8^��?5m�t��Z�K~W���)��8_��Gd[�7XD}�]X���~(��YV��c�����KN�8���^�#�е�r	Xۊ�n�	���0&�i]IŻ�fi5��rgd�$x� ������7����,��=<��7Ե�pzͻp��E�û��^��|S¡����\06����p����{�������ma�tq;';��O�K�2�.�Y6�hP 	�����v}���!�u/u����YG	�GK�(t]�̥"��UKg$܈ɮ���y���cA��u�{;�0�j�.�Ge݇T~��DH ��oVU��"j��v��g,pH9A�Ė���c�d,�o>)=���F���bIҞy�QW�ө�C��jvGd�2E�sJ.B�R�fu�t�Ϧ�'�sڱMr��`��S���ݑ�Ё�*��%��Y`�\	�`S�p,s�z��^��@
g|��S�r����u�;�N�i\!�G*����n�:��e�����'i=G�k�Žo��$vN��F� \���J)Ζ��̷-��g�񮙳L����~�("U��Y,Qgl�9I���:��`!Gvt�!R�lb�������;mV |��b��bƭ6��5啬A�4�X�e1[�Qcbg�g���,jcC��T���m�!�V��-�C������rc��5	���<��V8�ZI�D>��/'��bu���s~����Ƀ���}��Q A@����_ԙ�������q�Ϭ���-g�G\@��I�o'���Ъ�lm�m�ʘ��;aӳ�����:�<ۙߥb.%�G�2��]�h��)���`�1E�p'�D����h���J�}1R c��r���?^��߇Y�\[m�ղY b�u����ۧYY��Ը�Y� �%ϚN������o�4VD�n�}A��I�K�|vR�Q��oV/-�L�s!�5��EH��v��S*VR�%�D���.-�E��G�.����)�
�䎨S�g���
H�Us4�c	�ܲL���q� 3"?�.��O�Ԍ��g����V
�5�#�"sŒ&�-�}u�XK��ҭu�9jc��'b�4��ҥEd��n4P~k��4ٶ取t_��GK@�Z-��H�Sݏ�`��J��K!-���w���u5}��[�J�s�SS�&�c�]
>z�������s��ɀ��:�ޮ���g�%o�"Ð��1������D�G��(]����YU�s�'��3d@�Ӊ+GI*T�����r
ĳ=�@�o�[�o��U'z%0󺞘�����\���{�1���6`
��cFi��B��0ף=���~��Р�}+�<4�Wa/X
!��	�z���f����!��2���Uq&K3c^�kKq �}�ߖ&X��H�}7� 졕��
�v���*}�����_��{z�JY*7�m����ԩ�\����25X�G��\L�=YGT^q������W'�q�7K�6��nL��܋db��8��#2M��^M�o���k�ۯ�,��	nP��6<��19q4t�Ƽ\*;�Γ��5�I��uȓVk���Ѱ�
�hȸj�s�}�*�cY�b����VTE��\���dm����i5����X�1Li�5V��۩QiW���7�d���D�R{f��!]�=�WQ�l��3J����7����P��ן�$��[�s���aݢ��<N�6���E���8���<��4R��:5�����1�`�UmQ�w�F�N?c���&v����=%,jo�TCq��$y�M�j.���M(�N�!Sx'�c
� Hxd��(����5�[�%V�n��d��	۠+�*�UJ�m�6�\j���Ws|�O
�.<��/�rZ�H�Hp��ؘh�������#��`u�T\nӘ#���{���P�^�m~���Rn��c;�q�l0m������ԯM���g��}E
&V�=��ZV�p�_����)B`�t���
1�nI�J8���H��Y�_a?𑂱�.��b" x^b�E�9|�M�e �x�F�p2;Mt,$�_�i&5q��.��=����v�l�=�&��E���0-B�!���`�z��V�q	�7�2q��È�l[�CET���A�����Xܮ��V��.�/��#筞����(+����I�yO�T��Ҍu���&�rKW��V�O�)#ZIN����ꌰE��B9�_ݦ4��]��^��^$}������z�Ƨ� CT�����{�����gbcd�gF-���y�:�l�)T�%�u*���q�(Z�f���=�I?C�n���Ԑ?��$b)F�LUȮ�O,mm�/У:Ȅ:�Ö#�s7�3��_���!HN-�Ʒ��\�e���?��"s?S�E�(٢T�n��k��;�F�� �'jb�Q�Q��<һG��B�p�+��mǇv@�� ���(ۺ��Wr�';)���~7�E�c��%p�SɺnՆ�B���y^@w���>�?�@��*�n���G?�s6��g�A3�c9%ю�4*U�z�3
&��ʯ'4�	g�j�W�JC�~��ڼM�B�ꪋM[Ifs8�g���&���d9�\!���ױ���A��x����]��z����ӭՋ�%c�ɾB��� �S|C��F�b�+��2�;?�C�iK�8���Ż�N��{ή��	u,�b�I1���LhK씁U2Ccu�a��|�dJ,#
�C0��R� �pg"X�G�M���	�1����6Ky+�Ŷ�mΏ�	dgsȪ)�'D>h����wʏ�����`f��HG1��,���W5��<��H^wlY��eɪ-�<��0o5|@�]�]�蹄�gdM�W'�Ld��<6��|�*�XBߤ��2>���8�� �%����y�\����P�~f�í����gG�6佢}�X��G��k��F��;L��YA{jh�<F~�J0�g�:���J�~�2�%�mV���/����Z�,v��5�n5���l8h�X[@�αc������n�n.�89����%n[��J.�v"[�j��igS]���Xl�9p����31�)�R�dv�nX��?&6�"K����#�^��-��z�^����s�aL���寫������5Y؎1p��ī���X|�����h���=��Zf_�����a��Ǔ��hjK����_�	q�닔�g>B6�j�
��z�H��� ���\�&�N8��+Cx��T<b{	�H�q*��.%֊Li�������O���`�o)�p
LB��Kؽ|/��\��Ovx;J��oP��,?�'�,N��ý�5�����~Ï���yJ�6��7�>�*���ا��Dӱ��s�9��ܒ�1��Y0rd����6$�����C~��f]�Z+�f�2l{ꗣC�e���5Hl���ޯ��j���Z�+O���Y�J��b ���¾�~�|���PC[n�8��3 Y�_3��V���=g�b�� P<��	��x�EKFW�@`�d�l�f�+�-����S�yIA��j��0H�D$���X�V���g�C� ��|i���c�7s+�;��\���[� ��#��xf���@!�%�v�e"eޭ���
�k3e Z�!DN�	_CN�!�TH����oK{Q_��G	4��Bm~���֑��/�*�GY��ZR�aۆGe�B(��K��c)����neIR�s.� 6F��<�=�|�.���N�1��8�a�-�M.��r�ѵ�!��W���=�d*��е���Ԧ'Ұ[h1@�ƃ�̋�P��J7�^8����XsF�rw��!@E/�����8��2)]d7�^5���G%f�K��[��g��X��'^6.T
뉗� �Z>�v|6�-��̢��o[\y�X��h��vDB�9�ME'�+�B�٘�x���s@��+�2����l�\��x�X	���}2E�.���i18ל�Z�����Y�J.������uL!��������,i9�d^��ۃ�c^�z����T�[�c�{!�t��W<79݋NԔ14�#ڔ��ܜ&�#~�S�p+��P�������$�剜���<�����~�Q�G�b�<��&�w�ש��k�������#�������S�����.���Ӭ�T��ެ���Ѓz�<�=�I�S�' �-��LR^��������ͧU�?�I�=c�gw��cJSWwJe**����Ģ�\h�eőg+s�Q�1'����W���©���XQ�#.�Z�in2Q�	N_;?.tJ²��d�ǹۤ�6К�Y�g:�ͤ�(�y��{�k����a(��A�O=�)��'P��@�)��� �	��8E����Q��J]!EN3�w���T�!��aQ`���4NБ�i�v�g+�������c�9����3E%_d_�:K;����m�'l҇�R��h.xr|��jP�yUR?�e�x����H ��Y\w��F�2H������kT�KT^;����"e�x���s�,lC��ח@Z����F�}�LA��m�ق�������\BOԬW�Sز/��9?�;;KȜ?~l�'Z:�-���`�E�8�a���'a�����ixw���z�5z,�ww�L&���ZmK3��}
�H4��fcls�J"n��	`�P�	=��jx�_̒,�G7-�(��~4G.��$l�����F��A�V�=v�P�hˌ4���4��� ����X���^M�MRJ��×h�f{�&=�]H����+dw-N.��D��&�X�P���f����S��74�c,@�SvPV<���WT���o����'WKP�#�� s��zR��='�
p�mLl�y:>��W˸���B����]���?���g�jK�W6?�� }f��IϟƢ�M�>��Q�2��4NH��
Ԟu-���dk��%�Ž�(�@�Y�0�W���5d�UK����/#?¦�$��:�h�B٠4��0�{�$ѧIT��#K,w��*���:�W��B),-����]�p_@
3,n�C)�?�AD,���r?�hb������,@ɝZ�-�|��3W"�x@(7��OT�7/(�q�Gђv�f�s�,�i!	�k{���ܲK�H6a�k��B�xYz��4�?��g�.�Z��Ͳ_�L1�� C�F�_cM��\�`Ai8�_8m���U]I����s������w~*�J�ؾY��v��<B��3N��������mP*SF]��m'f�͆�ʫ=����ֶX�Dcytg��ٝG�iG��/���MH��1��L�P�V��Me�{RS(��|(����T�������!P2L�D#���I&B��X���k�ɓ�.���o��]ą�V�y��ۚ�"6�B�wˍ�1�^'�C��3�� A�~n�.-�=)��pK���5����+��u�u�E����p�ۜH��s��U>�)ܲ����EA�����]f�&5���GS���Q�lJx��qR�P�(+�]����+�W��e�x��O���Ґ4�2�+�ǭcf&�U�0R�۽q�,�2�w�OQ��dL�9�"��㈥tQ^د�V�n))�@	C�|i�U�����yY��!��_�0�[0c^"0xm�6م5�d,�|����bk����ȕv@s3,F�sA�\�1_�&��̪(���Rs@�_��%�?�H
�>���d���v�1����iƺg�l���&�Y޶��~�D�@���g���?G������S,]�4>z��Y��v�~z�k�V�u� �r������c7�`�hҹ���Ƈ՝8�`�d�����EVW�p�:�� BŔ�롗@�4�f��!�f
�"��r���|��^���� |��!=~�Y�oV*id�p� e��L4?���+�:'Vj�~��h�<�HE��^A���(��G�d���_�!�#�~�|n�6��� NȧL�{�ps2�=.���qýe�\Y&����_��K"�1��b��2�����!��|C� %��\ �����t'�)�\�b=��2�DWt9��_ �7��T��p�?w���8WN`pVb��)�Y�y����`}}@AE���H����H�P��C�T�\(ۖH�~�&D�RPQ+��Bi�	̻��>x��H�HmC��i��L�+�[$��N��)8<8���yjd���8%m��;�	�eZ
2�t�=U8�A$x���=��:������sUu����E��R?	fe������[0���H|�)�m�^�j��I&ϻ���ޑ���܋d�/`���x��舢�8�þ��h-ҭ���p;��O/�O(	}HT=�����YY�uT�R�Z��T\�@iD��W���ߌ焮V���߮�l������Ğ���`�E}���)nW�Q�l�Ϙ���}���R%U�U/���'���w�W Q�-�!j��M)�ǗP��%ϛx-H0
|E����@������q��j�(~57Z�^���Cx���X6G�� j+�n:}KPtoU;��;�����>����Ͽ$�n�׻;�WLb��@��M�!S�.w���a|E�0��F����J��>�������\�?�Nbn'��<�W"�$HH�M�{0��Rq�V���AP������T��.Wmu,S(_�2V_�Aw�꣄d�E��\�2��9s�(r�u禾\m��U����kL���]��(u�wG�v��÷�"H���3�H��y3�)�����c�-ye�oeG�r"D.]]`"W������O�5
�(֫�P��7���NO� �5����ض�j��8�[��F�V�"cC�8s�����U�9~�1�Ѣ����&��}�L���Q�i!�v��6��/�v��G��mj�92]Y�B0��YP�Y^:��K��ej�3��2#���Xٿ1�`,��j��4߮5��N�&�agY��V٘�H��Ą?��퀞�U*� �Y�(�f��nL�����,CS�\o6�"u`���\֪S5�Jo1�':�>D0�/��օ�Je�Q���F�B�@.1̾�"(��
m!O�ݑ���>Ӯ���c=��������M�ū_ORu�#�y��0�.��g�4�#�
7��o�$O8|6�?�)��g�F�y��;�P�)D+m�bR����ĉ��V{=Z^����@�f�k���D�g��@c��%�,Ժ@I���m��=x��]�|��IH�V[���9  �\n�Xy�F�	b�3�.�v.�i� �آ�u-u����d�:g�\|�\JRՉ~�Dw�ʜ���	���::T%�*ݣ1�=�����2�U��1Ү�éf��ɋ�>ʹ"L������B""[2�2|��M!�n��-]ů�]�r<FN�p$~I���۝8�lӅ��Y�m}�q��r�NV��1��v�>�ݿ.0^��١�J�AJ�3{�ۉ�w������]7j_ӿ�q���9��7mbo���BRI��q�6&<^�3�$�	�KR:�hE�Rs�۹I�g���&�ٲ�����@�9o�����Z��KuZ�'��3����M�տ�!���p�/�u��5��E�Ź�L��2�g�+AcK���ݘ@fX�S4�zkm���1x9k�8ąP$E���~�!��Nx���یBɏ���ڨ�����	� *����yC����R;�2�/�h��/p���3��ɪ���۝�+H �O7u8�
	Xz5���D�o����i��)�%Kk��m�=2�l�j��p^�dF�Y\����V���?�H.♕v4�K(�U۟��t�Yj�2��9'"G��$2�Q ����?�y���4N�b��q��zaËsH��f5���
�U�n��/��w�J�)O�Ң)�T�Q�!;��	G@���&̐�~ݴ�a
�eg�дf��!R��Ǭ�6-{�u�c���?h�xCp#'��2AW�F�����$X<�'_��2Û'�ޮ�2�R�����dc/�{.��� ��Y���űg�5dH��(-�$+|`��6�M�y��7��p~�n��Y�I��s�w7�΅�U�^���
�I��.�!�5K�ƻo�6��<}Ok����On<�I�G>��~+�`t�p}�����V�t��gO&���\֏8n�댱B���U���:[�~i�r��v��U�e�{��)�1��
3�KB��,xgOc���&2d3��������]w4	�6��5]��4�u/��QJp&@(�d��1X��IfsBf��
Rjp��ꨬ�4�|<-P�C����;쑘F��E���T�j�b���D�\X��	��m�T��n&�B��ޛ��Ø�q;@>���ِF�@Q£D�[ѹי��๐��Վ�%%�G�줸|�v9W�O��Y0����y��e��0eef�N��y숈S���9Q�a�ѽ�q�e����Sh�1�E����@�
�'�[�w��%���	�t��@�U��VoJ��	�$s��bݯ$�i�K���KX��1?�*Y ٗa�d�W0n�*01o�pX�g��DR{��S��m������<�~�����!�"����hФ]�Q��.+ː��%&Y�,��<�����A�h�l�o]�EśV}��#�@����<�[00Z�a�.�:N��������L#2Ԫ�j(o��!R���m��.�Ɨ�֋N֐H�|?���U!C:c�`��3/ղ�>��e�a�\��-`J���=�+�|u��p� ���+�#P5n��*n�g*��m�S��ƛ	�Ϭ�
�ߡ�N/�O�
0Lw�1O�N-�u�p�u��Ƿ׏y��k�T]L���%����n�t ���k1�J͸���C�I��j}K��B�H$X�:�!}0����;d4{P0�+���c�-9�w�6a��A$��%N�&�Ӈ��)�OF��t��'��wK��^#�2�S�P٥k��`�X�6d�A��Vj5�2˓�m�
�ګ��9������ad�-D�?��~2��Kjv�vb��u�crPf0�<f��.�w��?7
��u� �n/��l�&�}�mv����iq���n�5;�0�V�r�;c,k!�d��gyMc���@aǎ�.]N�;�4�V��)��N����Р!	E�r��0�"	 !>���h2�1�5~��ۃՐ��ކ�9Cw�}V��h3Ѡ��V���Z7RE�����߈�� 	�،tXV"Z'l�l
ӕ�^��XE����߂g�֫�l:u{�a�X*��rn�|��v�j��n!���L��m�pO�	�}��s�)��o��x�&�'�\LS`{��ӵ �����v]�_n��G���tj^�|m�V���^���So��`�@�Z$��+�ɪ�2��q�r9�t��l�k�dcg��L^[q��,�}���TdN%�%/W��SdAH��t�bs;o^cX��Y9��"J���y<����6tf��E��b��6 {�,�`d+�$7�C�,�B�=/�LE����6��o;��˟ĩP �d?-�an����>�_�T�iʢ�x�S�ąM�-���eh���^x]��{c8�e�~��{n��7!���������Y�k=Qu&�󰑜r���\��."X�?�M��\|ȮMrj��S�����9�q{]�������h���.�A��0�9%X��N����o�O�K��T�$��C��8?������C4�����Ƶ�}q/ fE�m��a֛dٟ�A���lɔ�X+dvGF޽�Ňe�Ji[m"�.�$�m�Tz�s<Ȓ�o����!+�ߚJ�n7�$�k�#����p;�13�̎�p�B}*�d����?��U��]��=seM��:KP�n�
x��)��j�TY�4H߽�"3��6��h�F��sv9�M��Gv#�qu�;M�^�b�������� "���A����$�r+	O�J��Bo�t����f�L/�m�FtLש��%U�(�.k�ᶲD����� V��;�2�n�A�����$�)Q�=-�L��򅓌O�϶�b\R��FS��~�Ǎ��ħ�����|�m�`��\*[�G	tj�.�D0��nȀ�������*������o9�8�Ī�Aq5u�?���㙅928�p�=n�m��Ł>=�P�JG&U�Y��D��qq!rC���x0-�e�xhe���Yh�d�<��6^�����%���:o{�k:�����s�2TS{m���.�g�<�J�Q��=��9KY�3^�8�gM�|rlR�����t�o�W�hõ�ų�a:/�9"��8A�``j�'�_A��:�t�"F���̨:3�YBL���C�?H��[���<���j��_��S &
�݁i	�Ƞ�Eb�����J�l�ýR^�}c��N7aV��mKL��>^bVy�6�S�N����-!�y)���G9[�Cw�N��V9�@������7,B�_S������A\8�'�V�In=��;u�_���k��*߉�%���_P�J�iE�t�G�J��w�[n3l�,��c���ҧ��7'
��s�������~����!М�C���u(}�f�y'%1�Ʃ:LNz`4�3�#��fp��?�9r�����̧��s5d��0�2�+ArH�m9������z��	��@H�X#��
�mM"���:	�c�/��C_���X?t�����-w%�l/�!₢��T�q����o/������hdȯ�����#3�_�Z/=f'��Z��J f@w�x��P�E�w䫞MZ��l�;ibF���u����϶ű�4OVSS�9a�`s�����c�J�9W�Bo�Ig�{��G�feY[+��`�����e �O�WnQ1B@��E����O���P�,�I��%x��f}ZW�W�ߐgF�S�����!~��ٴ���
�a#[���+O�=�Bk����eNν�	;6�L�M���^w��\�ӛo�ܗ7�����M����UY$G�Q�J�0�|(��.����<������k���K��D:��_'t���Ц�'t��D�K�SR������	N��1��
��i����A�r��߂�b�Kʆ�;Wx\������"tn9����~C�Y�t��8ڣiy������[��œD"��͙q@���s.�!H�^��I'�r��l�NE��I�)��������VFk���V� �R4.{��6
3:jjO�)�<���@�c}�tm��p,��t��}WS�u9�S@%��6�է:F��\�zKQ��1�LXĆ�	����6Q��ێ H�M7���bේ�Ȃ�:;R�ú����,��&�}PO����f��en�LȊPە���d�DI�@M�8:�q�/՞��{��s`9#_*�6�<}譙�dB�\���5� F��F~}۷�v��cpU��.:~����Krm5Ѧ�7��8�Z�ʥ�ͨI/�a�G�j�U�>n��j6�v�J� ��<��v[�����L(t1�05��ҭ��k�cy�aW[v����:/Mk`T�ڲ���"?f�m���^TYt�na�����( T<TG�'^�׬|�2��gt��d���q�dw�&���H��{§�]�N�Ci�qXlT ,�������0	��G�梓v��z������5�0㌥f2}��@ّ���Ҷϭ��6�`21��MT ��誰mt-�w����4�GgD8Z��X��2Y�C\ߎ��	�0��(v�8O�n@| axt%i�������VZ&��jcőޙą�Zh�b��Ɯ�l���(�~C�TKq�=���3*��N��AH��!�?��c�H������@ֻҚ+]q��>p�c����R'N�PU{0�"�-�,�MOw#��R��E����e�� ��yVn��&�K]*�K��H��ek��a��S���p����r��_4��"*�R6�>w_L�N. ;"I&
�����C�:N�D`a"\b�`�u2 G0��A�K�	wG�-�p��F3��l*c�	�2�Ff>f��*�&����i��&����$�3����K�1�>�u�	�2�TV;�	+*|\o'˞�(Ԃ�ÀS����
ٺ-#V $K���(j�-Y��Tر�-C�N���� @{_�@���>y�A���'S����S!M^[�v�29�\kvJ��C��Dr_����F��3�A���;��AX��V�C�F+q�]	atB��;-C��>i��k/�}e�M�q�X��M����W�A��O�?^����N�=.�,�8V�6鱂7w��c[�͛󚘠"��Æ�+�Q�d��Z>HK�&o�aIKZz�oE�sp����-�c�4�{"_"��e��RGu+@��]=�&Iw�8Ҋ(��2���Ș|0aF֛P���g}+�ę��[ș�3!5��4XU?�T\���R}�_�Y+�o[&��@d|kO�G��8��L�{�~� ����>��_u!F̴F�Bo;f&S��ZQ������[�D�L�D�l8����y����8n�"�������9U��l�EQ�K-��t��	;�@q���� a-wA��y"�f�cT�h�J��Ȭ�f4������3����� ������\�u1X���Po?2�Dۍ�w^f�S�Z7�S�o��,�L��l��%_H�� �6�u�'A��^���F��St1(��_/�YxrS��i�Wc{F"��G��^2S��Dv]�>�4 ��gaJ�US����N-���d�&C�HCPF$x褨
i6�i��t��UC�-xI(���})�0�xwwD�ux+��,��u2�z p{P��Pg�撘�\��y(b[��`}�=d����$l@�:J���)��/�H��,�O��c�K��&�fc
"�gݷ���xa�TbZ�nJ�s�=�}`��pw��%�pY�uo�|	^G�␕��=Pa0��;4؝��'�4{ 鞰���f\���X�Ĳ>�^���q�1�0�(oLWW���X~��o��wD3�}t!�%�����vL=Ե����M��t�R�L��^S��j/OO(�8ƾE���t`՗IPDc'rB��b�_a�qXϳ�[>HeXɰ�t<ޅ.�a�C�RJS>v4%��w\�2h�l{\��KQ�����U��*
����h��4���#�B�Z�(*#*?����>=��B%�<�k��J#n}��O3������ <��sZ,�U�&���)3���g�`e�/���D��?�l�&f��K`CA�[T,�o�~*��� ��� ��K3�W% ��pO#(�2Q`r9�"ӿ��J=�V�q]`	�/����.f���J�@�~����\r��n.eՑ�z��2�Y)(3E@��l��{XtP�Rt��x��ù����Ү�޻'�,u��p��c N¤��ƺ6���W��P����fԽ /SP>S�����#2�
�^�=υ*
�zA�Q{�oy�(��|�X�7o��R��&�����'�0QXV]���q��u�F8R����3��IV7��!�9gi�q�ͳ�� ^�"��#7�)��|�^'��'\��o(
j�7͍Ǻ�<`�.���KQ�� �Ѭ~�xsE�k)FL��w>�� ��X*��^�o�AȎE%�Ms1%P_&Ǫ;��C���9:ah��-�[�R=��4\Ɛל	�JܛQ��y0[�:�΄���(O�ʂ!�A�8چ�i�|��~wDz�`�14[}	ʴ��&j��6�y��|E8Ό<�"
}�1�M����$��0B���=����AD�hm�d�;��s�k�2�|*k�2�^?0�!K;%����<�CU����[_�rn5��5���;�p�Ӎ���))m�N}vGap��#75 �6��]�:��)"�����M�E��vV����Kf0<���&�+K�����^k�4=e����
�9X��:B�R��X��Y^��a���l1�V�������C�k&��%&�2Þi6F�cDQ��d�ם�f�p�C+���2�������8�+)#��Gfj~��# ��r�D�G��f-G*ٝDװ�Q΁Py pup�@��s��� �y�z�Xja�"�\��6�i#��ھ�"��M�����3Z�E-�a�V�9B> ��DݚgJ�$�ʭ�ѝ��^4���tė�!6p�e�JH���e" �R�$��V$7a�<�'�1�ᜅ�uӐ>�2���y��A�S�Wy�n�6�0�凾��/��藤$��'�%6�6�P>��^�
(��Բ�";��Z���ڡ��?�L#h�!4+ �;v�NSs�W�����7��k��t�:z��6�]���t�B�@��~��6��h*ӻv�[.�f�ߠ��S��
�������Ǔ��7zA�{g�=s�N��V$F�]>�2?Bhσ+m��M�7�Z��֢�"(.��wj�"&����4Q�,����"���Q�u��,��\��*XF����.�&��4����G7���?���w�}�C?0=��n_܍5M���}���dT�0ߕv��FU{g�c8�!pH�d�O�F���q�k�B����y����6�*�~%P�ί5 �J\�]����mw��G{�#t�x+P@�KOX�3�b"m����^��N�rhW�g��c�eq��@��X�+����՗�M�v��._2�M�}� K��f�IX=� �d)/�
4�yԔ�]�et��Wт�#�G��_�����[��1.�8`"�I����ɵx�xbC��"�w��Mҙ��7�����9W��uZD��u��K�M�
��Z[q� ��m�j�(�gZ�ES� )W4#�l�1ds0��\���`[�c������Omڔ�.��.���b<��0����#�����dЗ�r�'w�l��`���03R�5/va]S���ì���{Ҳ���m��*���vB���c]���8;��o�s�wo��֔1=�1o]���۴��!��[�j�Z2���-��!>�}%x֣H��Z�}�|p�&�Ke1#�tQe�î���c{b��Os��ކ��x�0
��p([�|ATFfN���l!$lw�f���{'��UW��5�o���Lo��Я8:J$��Z���� �����D1֠�(e�ˉO�G��'�_4mN�*#�(pK�p�7NVu��:$��m+O�����:�)�FO`�{���t+yU^��y})L[>����p/��T���Z�]l� M�[���{�v�!�,�b�TR��r^��n�Gl'7��H�P��/��]]vC�3^�|ߝ���)��mܲ r���n� n�oUb2�6�=�x��Zm�a��?s��'�|�P�|1��QdH��ly������'�Бܧ�7~��ئ��#�Ɋ�	�� F���KűLy9��|XX���������2C����i!�t����6`���$�m=�1F?��+G�"T�q�+�4�ވ`.߷��t_r���L1�*�������.R�oj�`�<5����V���J�1�Ty�ws���� H|��Ľꃈ��V�j,�&!����h�Xp}�@6�O��
nA<���d@�+�l�̃�e47�7�s%��8���n! �(�*_��s>�R8��71#�k�s�m���d�#Ɲ�E�&�]Xg�j[����j�$2������
>�y<�	ss�<�C��HRm`�>.	#��u�;���%��{����R���`�;���ʧ��6��y@�� �d�Z���� ��x�N��B�⒰�tI,�p"���t�y�B�&���I�.�0�+�-��F�ߓ��%�8U��j����6F(�����i�T2����F(&�R؝��3��hO�@C�i)+_A3��O4T��NBx^?@^�iR�q({zP�z�XF�g�F�eE���󓞥,lXW{�$���S��\�� �0�K�*� <�
|�
������h;����(���FF�O(���J�+��:V�74,��|�)�@7�NUq��p¹��C�hR���y)�R�� ���ؓ�E���ܚ��	�Τ��T�G���2�m�""�,g�����j���뛖��4��`% M��iv�e�P)���j���o�	e�"�2�cg�ݚ�V.>�����ej��o$Gχ-��Oג|-Osn%�ͩi%�ʥ�-GfS��>��y
	C�lj��� �P�I���� �� R�	��%w���;�	�#k�ע�-4�����ӿey��
������r䕄4��?(FQD9��,��$�r8 b�������(�<	o���>��\{���O���� A!����-�菔'3��JP��Bǅ�J��yЉ�������0vTr�3$����6n`�q����-0�'�t�]pY
���l��.��C��wi~�P95��r*߲���%z	
��%C�=�~޻i㰈�"��<ΥM�������5> @�F��|]��b4MN���e��w�3�gxp���Li˳�<N�)i��]��"1��R�����+xs��B �4���;���S���|��f�,������~�8^G���Ғ�����D��,��3�޾��3m[�4�\(�r 
��m�_5��u0O�*9W%I�U&����2}�0�w��CS��w���م�vCؖ]�*��Z�Iۨ���b��EҖW�8��hސ`\�����ӱ�w.�%�_���c�è�OQY�_7 n:K��?�G|"f�t�l��-�c�[7*����؝~S*ɭP�Τ���rW��˫{�1��*���([�:�ՏE�0z��sl�w�r��&o��1��̀l'������V���7Yd��/wU}�����j�B�mv��dS4�}(7��?���ߧJ{�@�j~�f<���� �F�)J�
M+Sf�?g�El����{8�@Y���V���	�B��3��ܲ�XJ��-�~��J���'�w.��!��o-8��d/�C���x�@1� ���c�D �wa���1�_��uX�"؟��ڲ��h7t?{|�{%��Cq�䬽z��b@��6yx3Ee�+�@�g	�m(�v�҉ޓ�ێH�������=����[�:�vF�v>�K�J�b�=����	�Ҟ�Tz7Ƅ��A9�u�ģI�0�����qkY�&�B��Tq���q4�h�cө5ޥ���� $�ୗ��9O����k�0�Ul5@����de\:�Bu.�:��S��$��S3�����Q�5�>�,7uoQu��$��C�zx�Ƅq\�Hi<S���4�`�x35���s*�}��(�v�ާ��C��h�O�JA�LE�������Iq���ma/O�nN�*/[���ai� ˸֔>3�L�40�WWB�(�Xr�;�YVd7���&��N�i�Ԟd/�)N��
��Ec_�}��ZW8]�%{��y��%>�Vk� i#��¦˰Z�z^J��>��v;�r��L����!((���J/�u��.�&	!�mJa�����d*����C+Mܶ�)�h��:� �'������iU����LU��c��7�d ���>�.�j0z}^ҁ÷�����������w0m�����m�R�Ӽ4�v'�cj�?�G0�ay��/OtoClv'�,�P���$Y2��Zs`�<ã��o��B��h����3w��6>��,�5R�.*V��k/[� @�ܜ����u
�{/x�Kɩ?�!��v���ܢ�S
k�>�Y봅����E拞�J��)>��b4��R#�j�#�p�I㴄Z���p@�r�� �WQ^�P���S��*M�ԇI�>Y��P�!��W�Y^p�U r�(Ȗ�^��PAY�DB���q��>V������I���$r��j���2qb�G2�Z��<'�f����(�j�V|p3��@+�{+E:��ʭ�v�G1��$��գ�B�>�%L��t�B�lo�g����tH��S$V.X.bƍr2�;qA�y<�:}���oƉ�!���j�7U�\HC�?S�uI��M/�M�sӜ>�8��Ag���F����oJ��^=��������N(�
��uk����Uf ���̱� ���u�༿�f^e��yT�
I���ѻ�m�}Bv��s6�UTlq3�ga�uxxa�</3��6��H��rS ����Ҝd?��ΝW���;/)�K�� C�o�����Gi�4L���c�����;����7��������Szdq��̓;cM[DD�$�eJ�^	 ��FE]���vbG�Qٲ�k�P-ѶX/��᤮���KІ�!"�Rce@ ���d�jÕ\�B����吨�:/:�~0fA1�sRt�>`�s��T1�ԆT�v�� �.�H���l�d�٪��:f�6����IK������D��y��L�N�����E������,�ǥcBwQ�ч'�)�(�ǩ}֘�S��vQ�w�ѝy}4�P�ð�QŘ�b��5�rD���2$��ʌ��˕$ �pŊ"=�ĳ,���m0��kӶL0�t2v���9��8��hR��#���&Y&�&��q�<p��=|O3I%��p��	<M��˯d��r��^C��i�*��%e'� q�r|���(_Dq65���ԏ	�k�zM�q�����W�IG;��Idgl=�\��HQ]�o�����j5�P����`��왔0˟h��;Ao�V�	���(v�_|<��IնL@�)n$/���\�����˩0Ղ�H�	l�>���R�������;| �4�^<��Ls�3`�cq0�����@�zIZ�������d¶�⼎��[�ŝU�˨+[���ϐ�'͗�S���S�%`.fe锇S�����>$��"J�螷�~�v����gt�YN�1x�+�_��:g�a�܅:��Wgs�.��)fT)�� ������rj�A����|%���|�s�#E���"$�5G��C
��\������\��a��^6����,�<�KC�I�4���{7Y���b�<0�;��ZF��!$�/��4lT�s5�R&o'�`^7ysDY$����f����)g�0�������GWHh���ׅ碳�5�^��]x�Li�d�h.�9�Qn��[����1��������rK���������ka<�u9��T���x��h@)k�H��ڣV)���z�A�굽��v�yc����e4Qݝq�1Q q�t[���Zm�^��	Ο���r����������U�7�����_�}���`Q�r7��?��[¬P��	?H)�q O�|�pK����B�fW;�/au�J��U����Uc��]s��+�C�#G;eq��O�.Zrk8��_�9ĝ"��m�@�4Y��=��M�yTѾI?o�_�F���Ֆ{����`��2SY�$޻M,�����#L�{V� ʏ���g[��
�^�È���k�8a@����QH�񐶼�=�!�˔��Z�
��mGClL�c`;-H�j�$���ŀm<�[��g�����Z�����ωH��3c�0�<"T[��j2�Q#'��(��ڑ�n�5���:/X�MC"�aaC^]��F�]�W����#�	����4���v*;ST�e�1����X�qgL*��VE�-Z�G3����ۮfT�e�]����N6yT��*MC�����u��-��iU�����"�֣��/�1p���2�GAg�z��q�]��֚A��|���:��龸��f�-�%����d'�[Ģ�`5�Z~����X$��^�}��y���_��p�h["�G��3�#�N_�G�#�n_�y�·N�0l��'�2MF��?b������37�n������cS�N����
>���ᖪ��}X��dOI�����tt�.��)��mr�xF��r�Ĩ�Ն}a�IA��9Vk����s_�͛�E�D���,���|�k�ȬY�w�X��8as�:T��}�9�ΜY�:E1ˈP7�L;���JZ��u�P�'xI��{�o/H���1_"�.��a�9v��^�i}�~�_��k���NA�s�������?�_;�9K���*���/8� ����2�}��G���X"��i�g�b���X��m�]oC6;9 8ٖ��Hn�����$���1j[�Mf�^�숧VS�'��R��JS/8�:����ϝ�F�!�Cd-�1a���a����(���⹽~��}C��tv���^E�"d���Cl3{'d�_���/��
Su��)�l.��p�1�31���������2��O:�%���ĳ�u����l�6X�3Q�Fm�θ'ؗ��j�*��"9�"�)J�Ռ@��O)�N�6"]uW@��]�o>M���gFY�E���o�\��W5�?e�FIB�\��mEh@�k+7������ӄP��h�����0QD��BD�|�
��)}{����Oݘ/�i�<�T]Ҵrr��e<��2z��jv�|�L ��i�PJ�Q�7;QP�����8K��aE�8�cL<R�!d���Ir� 
����ƥ��(�T�z��N���2�k���(�:��j��wh��MrV'�Q��������mO�įV�o�q�W��EG6�*>rx6_?��\钇wS�p��@?�]�2�{v� 6��5
���NA2�6كY��S\2uZHt�T>�T�z��rX�OSf`�4���}l3U2��Xw	��[���G��~�3y�:�#�Z���ev�n�y6w�+T�����Л�^� �il�lQ�ؽf���V�O‥�n��7�����W����Y�H��*�Ro��JX
�13�l��K��f�<d�ٯ��B��g�5�^f��*@�Hn<������qX�m�w�p�J��m�ܸV@ϝ'j���Jy ��N����Y6;�����t@H7�v;~m6�TS����׫Ԅk�,��� %�
[��a���z����h�wUe�oB+U�9����!XG�W�@䗜t������q.9L���CB��6e���Sԭ��$�����Tr�xW'}J����5` ����)q+�a�<*�D�<Z��=u�)Z����,�xx�G�1�]`�+p%�+�|�=�|Oj�Vi�Xy\�����C���	�=��L��o�u��`���t�r�F��,�0���:��go���:EC���z�]2K�]-��E3̕�� ^�b�X�is�e��4z�,���M¿��ܧ�Ds��) �P"���+���	�uX���Ү\3�}��7	op\���"�C�i��B��aY���A^��J3`iK*S���MΪC��f$�{Ǜ.�cF;������o��MK�g��wȘ�c��7�8*��<�U��̄�dd�C!ɒm�q��"Z�8?w&�>�C�<ڢ���P85�Ute=�d��Z�#GR,��ir$������H���I��'�v�j�Ϊ��U @��
N��=�FÏW��ckz��U4�"�t{U_څO��Fb��i���<���^-��q�E�N�L�R�7��0�8�Hٳ�B��JG�����AT���֦/���^�n��D��6%��[z��Ć@H-%w������������yˈl��n@�P�ӈg���"ѭap��X�}g����?#.���u.w�tt~�|�{c�1�Z�2W���v�6�þ�#R3�4�@�;��vuyX��糁>b�C�T<�w*ZZs�?���,��>��Tkfo -����w��ؐڹ��-qW�8�9��+���������濷g1y�%u�xZ�)=�T��$e!CN�\9l�{��p�s�m��t�˾�@�}���Zn�L�S��0�G��!���/rT�㚛cr�3�G�47e��]/ܱ��P"|g�"�M����'�\�O�ʯ�n�n=ݷ��,��܁��3��"+H�I
:�õ�#!����@�v���*��fdsV��!{<�<^�?a)8�ۿ�i��/���)�!=�8�E_�%�F�e�/��A�T���f�fE�C�?���ձ]0}��t滭z7jp�m *�l�.���K/�9����29���Id�j��W�#"G�s7�,��:��O�3;H��&�@Tډ}S3H�o�Y��=����z1�K�r�.{[���	���>LH������WXͻ���%s���Xic���YZ%T{$n�a1'���׺�z*ݴ|]_uX�_��t+Na!؏�>TG���qT�a����dt�!+ b� �_%u�����2���Ԁ �Vf}L�^K�-�� ������Zb_�GGx�Ś3��G��/"b�����!]����G�Y����5d��V :��V�Sk�n]ڣ]h{��l��C	
����6#z���&��o�E�, e��u﬋g�Aw�D���?Q���Ђ˭��?&S���N�X�3�_]� ]�$��pKj�?�xg���K�y>�nf�����Ƈ�qݎ���-�yc14:B��܁J@~\^���������K�4)"}�v��r7]�u��S�kx�霃�`�r��C�a��WeD}�6ژ�s����o���}B��2ז�S���?y���c7�S;��>�[�4\�|�s��;
KX"�:����n�Ni�U���WxI]��"lO�'q��v��E=������E�&j�=Ɲ2�-p��|F$�K��eo�o����}�>�|['��:]�TJ(;[�1[R��G2��hdh�./�o�3mL��A/���W�?U�8RinƦD����`���:}��B�� w.�@�4�����X|{�7R>zc�OYrP�TNQ�]��3���7m���ʪ�?��
�����6��f�P��_a�4��<#��}4�Ra^�\��,�����-�n�d�"��	*8�0��SY/�_�qw�YS7ȁ��
>��-bN�R�D��U^j�:�G�Y���B!Sdw�fƥ+tĲ��ּ�f�_�m��`�J��n���ϤuC��/�7��E
z�i��W�T"��v�y�H[��e�*%\�I&�?Ɯzؿ�K;N2ǐ�S���b�Z�w�����΅��aOI�ʗ��幕��]�-���g�d�K�� o�I��WPL�K1��,��}�@#K�FR)�R��D]���9���J0	����	U�W�^�4��z����S�0��0�u^B�	�1�l��6�$P���g�sؐ���iK����B�E&����g"1�m����D<�a�א��I�7-�����E�F2I��^��i�4V3��ӽEw����b�f�LN� ���;<��!���e����;�7j��>.��
B�kngR�9�-����a�W}GPB�06]a��VF���w7���17tn ��Mj x����E:�1|��W��(X%sm[������§�,�0,�s�QYi@u����h������ �KJ�w!�ys&7M�3������N����5����r3����S���d��''�/nyh��D�[��/���j@7�NMB��'�}|��Z������A-������v�ć���ǼdQ�D2b��b3W�i��>��!5�f�-$�-���2�1�Mi�����fM_k�B�� #�eXm�ON��_>Vm����z��_\)��)Hu?��bI��ʹd*�=�3m	%��H�����Y"�k��։���{��UK^4�d��3�il��D#�aN:���}a��d��Q(]˜�X#����i"lyA����ȸNw�/���S�a�u2��FtL4'�[����Lͬ�NS��r4\�M@�|%�������	P-���aR�*)�薹���eG���'��^������5��v�E�{s�ڴ�������H��y���.tM0�T�o�-?��/���b�49�,�5��{�����Uh����|)��d��-V��QvV������@C��-ؒJ0a�h;N��_����܆T���)Ӽ#�0�?]�����6�.��PE��x�I-�0���4:@�T!�X%jP�WP�IBgx�_H�ߊ��Y��jy�!����
GKI��[1���JZ��j��d^���u���U�dpU�0�N�=@�oN]�t�t��P ?�\3X�hѤ暾�،��ae�J��x�6�+��M�NG��>=ܱc�[M��욟Jjw-�>�'P���U+`H���S;����U���L�ǥ���vC	�e�MW�C�p��_cB�H�!��pk�ۅKb%�}�JI��D0R�؄C��)��9���f�3�59��B/��qi�"V��OIϙ�N)䍏��"�Kc��쳋�s����-���.k�-��(��0;����(��-1<��v���k!�G(����@���1y3�sZ�7�"n	�Ũ)3�!��x��g��/���p�!<���;x~O�}���ϑ�wk&>+V�@�o��Ķ�(�_���'+_���t���aKa�91�B�N�N�?��M�\��G�A�^f�KѶK�3�L�t4@��h�$�k�^~��-�߮��)���0eI����V#�U"��S�py��t���Z�8�h�Nq=U-�RH�Z���,��:��o�Y���e�@�d��[o�++�V_�R���	��i�X�r?Mt~���˄���d��+��cdd�V#]Q������� �X�9�!Y��� �|��!�-)�!��a�~oj�JH��=	�!n?��s�z��L7w�kó�2�V����18��:����_#\�$�m�SR�6w\-� �o�:����!����)���e�)v��\��-3�ZI���K1(�d|9%Q�//N$T�@dV�7�?!t�.p�(��8\��ת���T4�k�ТLb p��Z����j������/,$�Tk��������o���[�4/:�[�I.Brc��_e���.=Y۲ ��Q��7���%�G�3dF=A���Á
��$<C��\�`w�l�bi�����ӄx�k	A~E�Ԡ砲�Ei�MЗK��*H`o�S.8�<NF�Ѻ���5���o���SF������]��p782Έ"�N�otյ�l�/ 9�i�}�YU� l{�82F�ч`�Ɛ�F�k�#o<�ĵIG�u�Su���L�qP)���*����V��z/õӺ~��� �{| dD/�4��yR�T1�K96`��<h��'���5���5y��Yi��������H��n\쏪Չ��U���s@�Yy���9�N�Ë�v���3a��~�Y��C!LR*�|�N��<�S���9���C�=~r�ϟ|���q���E�!��V{�Q���=W'�{�~]�ki��0@8�W�m����<&-�~<4G �aM��羀�J�Q�kYR�S/���=ɖX�R������������`�b�y���i�__`���"�.�O�$u/w�g)�F�п@���m5C���0�A`E(�D�D��+�wQ�71Kh�Smňl,�nD�&P��~�����u�9	����=�,�j��L���0@~�(`�6%�'���KX��|�i;K�61���tl�1�&���G������B�.�f���wEr1�uvsʏ��|��qz��kHzE�@Y�6�&���D,T���u���1���+�d���_��;ƿ��Aq�q��R��¶6��ZY�-�m�$�T���x-�D싏8��;��1G��;��F w�L���A ���M�8���b߾Nbu˘BV�0���>S�'����R���9 ���%U�^h-{��[����So��g}��̹V��M[�L+eh!�yS�G���s�H�4�k�7 �x��Q�d���;��<O�;=e��I���2c�F(�f��1�m>Y�M8	[��n�1a�rt�(�U�'����n2��Ad��1z���U$��l�IY��I'�����ݣf����#�*��IB��+��P]��� J����y�{���+�t^/b�[�SR����lbL�Sі��d����8��y��)n�ӵ�Y���z��|��7M޳��`��%ԑ�C�>S4Z�g�I�2;.�9�������X�(cG%�T�9*�W�������X�����r�4��B$S~#�N�V!΍�ة����u:�K�N7��{=�¼����{2�`��UWcs����r B��J~i�����7�7Df6x�s�m��4<^;c�^ꤧ؏��{��	F��������\YTC��9w�+���M��Hhq������>(����e�0�{#;��9X�1c"lf�H�$%/�U�����;�EQI��[�q�5����T/���w�4��I��H��\Q&�����n��6����&ld����J�l��t�`ܼ�D�r�0�X��Lz+��H}%`Un��3y�/�^DbU��<���q}.6�U�/y�N"bV�o�'f��!L�t���)��ߋ��h'��k�߆5+�c�#���v_g��S��r�o�Ճ>d�����3zzfX�w�jIjcqA�ʈ�ʦ�sT�4�n���9�,�2��^�&sN>�R�C��J��0�\��������H��*R<�%�ͤ��|�Qt{>�A�4sc/xF�<�'=�aO�A:�u�_���D[�����V��'��,a��B���!��*�!?�\�������ϣX������;��|�ha� k���z[:>����|?�����U���"��1�7����8�O/�k����B؁��[Y�~Ӟ�����e��f�e�U�P �?k��mիG<}�'s�:��2��1�*����gkO�cFE
h����ŗ����7^����x�N���H��k�r��u�ݿ?����B�`�zT���>���r4���v�L�XW$Lb�b�ٻ�J��s:�Y�ԥ^�ҕ��l�9�rn��f����9�f�Z�d�:Ul�a��{X���A��=VtV�@H�
Q	�d��Z�0��o��D&�1Y� 0���������d�u�6ÕP��)�t�:��ꠕ��Sf�,s՗�_�%�6TS�qK�dl�Jo�O�c)B������a�6+F��x�����Z3L�=���i�����>�	Ԩ5S�9j���f��̽�K��,�ѯY��f��g�2D�������J{P��ө�-V�WA�׌]�_���N�[9���$<+gx8Dn�rt0�a��0E��z?�8�=+��b`��9�Ϣcu�'h�!��<��[o+��pW�n������>l]�t�8�v�'�ӝ� ��j�d���q�����(�p���s�.wjy;�_ɍ�s�&ٺ���ʬ��.�2�.����>1�:*�Q6%���U� 8A�+p�T{���ku��M����9��?$��jc�p�F�J��j6�i�z���]Lʤ�:Gm��T[,6!����C3y�7�
���~v;���@
� �j��e�h�ݓ�V�_R�e����@�+�W&��������y7&;�0���ⱒ=�ь�#B���̟ 7I=�\�u�@V()�[j�jlxV����6T����	�Ѹd(.Zl���r��kXJ�v��Q��w	BE�l񛤡�d����޾��ϋ��.ʬUEB
4J���]A��;[p�R�@�����0#�vcM�]��B��+'�t�t�t]ib?�o�Y�(���r��E+J�z�ʡ�9lj�:��k�Ҡ�=�W/y�?�$��[���SR-1pO%`%7O�B%i�A"��
	��5'➢Ӻ�$Ƅ1z_p����Ț�L�#Λ�
6q�%�{��&��7��o+�����_1ݨw@��P����>���d}���u�%�L��mMx�$��<Zf���@l��㮞�۰F}��ys`�+��<?R�@���C��Ƈ(�I5�a���(�)�$���}d<H�d�����*�
�d��#��1�C�Ȇ�݂��j__b6����B��I#�ȾF��I;��Y'���-��z^'���rô�'����s��dN}"L}�CW���"-W*�
�πS��PΒc�Y.���fl]4��3Gr�uC�K�,���Qm풏u������kw�����=�и2f�������\����VmU�����dqo����ĸ�A��͆�̂�0���<[�"p�Jl���6�S؂�X�D�|I����eaǣ?�X�LN��!ʾ呱��0����Ѫ:�ށ7���IvM~{�Ԭ��t~��1eye�7}�����߿��Inl�Y^̣'53�!u���ф �B1���B\8��cV�M����Cgj8���f0=�m�xV�&�3±V��Aҳ�w4Q
����5�@<"���=���<��r�z�.�).��J�`���-��tէ2��Խ�b��So�P3$�Nc�Z��-9[��9��:�Y���j��r�4���E�89�s��Y�����<"w$�Oi��D)m>����,���(H^-ȗPw�2|��3��&Wj��;�gX���L�s�����6�gG|������҇*J~�j�BHgX��Y_��0c�5����&������w�}F�/�M훉Mr����%�߳7���X��������TS�>:o���G�¥W*�Y�ر�r���6qvVөb���~~�>6�Z�,W������t�
��/es-L1���61>(��+�����~G�u;p�A�ze��D�#�BC�2ƭ��M�=�`��yV�	�W1<u���6��wM��<��༓���*�C����j��A�D��m�O&�8�v�=��O~ȉ57�veNvu�;��Vʖb~����
���� �J��#R����k�խ���� EC���|r�E�l�
/���B�]|j��l���%�$O1���IL�rer\�:E���NZ>7�~4���1Ծ�u��^Vv���I&<�����
ذ����P��=�6]H9*����)�Dy�Z+]�/Ƈ���]��f�/*fv��snk�0q^� 8�C�27l
|h�Xq��@���E9�#��������l�%^<�bjC�
�f|(T߭U���8����}�ϙ�j�8�C���v|8� &r�W:��mf�n�t�����1�� 3�2�{�^��&x.X9�Ih�e��fl�3�o��Z\����
"zQ��n��#<�4׺q��sC��Dk�>Y'�ѢN�(�G��U�wgj�D������q��ɀy�B����A�K�A��~0��Ț���}�����wM��c{!�n݆|��lqXp�\ڐ�K�R`)�m�V�B2�+�?J������� ����.�ce{s~QS�@T�w5�[���u˘\�Po^�������;��P���M�>3I�'����R�/a1�A����ݞ��?�W��=4�U���{Np�O�� �H8.��݋3��0G�M�{����;��}Ͻ���sA z���a��d�-�����3��mF]+Iꛕ��jOs7r��dc����ľ�����Rܧ��Ӷ��K�uP���|-dլd���|D#�5��@�X���!F0 ��ZQ��*(p.Or��V�V�v��ۏ��W�j��g���R#�Q��(E�iKW}S�([�����f]� ������	=C��0�W��{�)��)Ô
�(�JAOS��C���x�4�*�$ d�{���PBVz	�M �¡o�vB��cG�����w�.F�MM����r�&M���m��sa����_�o������g��݄5�|�i�%:��LOo�DO��0)݂�-�oLDm�2�Zf�:^v�np��Ix�Tv��1��4F�K$"K��"?Uw<���<�z�Y7���P�E"$�N�mw�^
�Ƒ
�Xpjh
�����b3Y��)z�O.Ӌ6-�e�I�s���uԲ���,�?�:X5f2H��ټ����0tgB��;� *������8�}m���b(�%�2F+Я�]c�~۟1E��";��&�cH�ZP�b##��yÅQ 9FG���4��6��X;$ۑ�i���嘮 ;h.���m�G�D(���[%ǻ���s�
,~8i!�-��()��!�⯜�<<B�eR%��"��?�7*$����4�W������-8����D��8ݾ@b�A�H3~s���MA� D��P/�Dx������ʖ�+MlS�A�N�aj:�E+����N�+Pq�QJ�/)ܸ�����qIJ�����V��%�����;;�Y�"�b�]��(�L�I����{{NJH��j��N*��+z]���3�*�V����C���<`^K�	1�Ʈ��d�/�0�L�G���ÿ�Z?���'�y@���B/⿫9�$V�K��Ǻ�{?3�rn�Z��0N%�r7ٱ���k�/|����>�1���Q�[nF+��ZVQr��1s�v���*`���"ʪ�Y?K*���a�_��Q���9	?F�Ȑ�T��]F�"�\`k�_�H=�퓏U��W%x�D�t�d�
kjG���J���a9�����U�O�!�u�G3�)�s)�Xq5��fݑ_��K���j9|K	%-g�� >�0A���蒖V��8�����z���r��G��:��]��g|ٸ�q�1���v��n"�3 y��n��A����'�h¥��	���L�U���p�#A˞�+XD�Pq,�Uz�ptYgo�k�%L
Қ�~O��@�X��?���׸�ɣ3��ÜqQ?�O�j��\��301$~����Z�(�=��Ꝏ�Q�X�>m�y�~N�j�W���\�*��W�w=�Y�����Q�ah��v��`�x��,�X�R�R�..���F�b&L��;}r0cz��E�(� w��?0a�ă#}�Ƣu�c�Z�o�Ԁ����x8�X�w0���K�a.{P(�*�h��˱�l$pCy���qv3���I>;܈�=��bIv���NQs�riМ�0�Ü!�+囉`PKx��;�U<�)Q���}�� ����)�R����g�#��H<d젒�����U�w�sیGUq �|���o���Y��-�k�f���/kx��?����`��^���*�����+��L+Ʊ}U������e/l�6�m�zu�aGP��e>kCnugF�lC��X��8�xVmr?��z]����b�m�ϯ��c=[�M,���'�pCR��a	F�U~����o�2.�'���@���~��E���9���w��!���%^�~�&p���#2{z�WO�]�M�	V�j�i���������0�ȥ��\ �a��Szu���v��*2���>��0�0+�9`р��@/a6%�Dܧ��B"*����Ãg;��r"q�|��|cp���ᐕ4��u�xf��w<��ـyL����p5o��1�����	]y�k���v�>���nK�M�8�F��X)���X�t�`�"�Z4}m^��+^��u皘d���8J�v�"T�F:�����iv�� �n%���r�e�kYrв
}3����1�~���l��;Ԣ�sJ(Fc�` >������=h��!"��ԓ�@�s8&/�z�5]-�0Ab%�����p�y�/�s�6B�P@ݔ�X�x|��OrlZmt�O��~�F���Pj�na
����i�ړ�թ�*Y�*��׮S�S�V%�8��"��6��hˤ�"�'$�=�).��ce�q�\,�W�����;�}h/�=��'6���@hpk+-�78ە�6�r�H�O���M�9��4���НMqm��A�ohc��l�B��*�|W��k'�o��k��A]T!�'5c�v�����Qv��ز.���M[+�K��c2G˒���ޟ\^yIi�=�৑��7��ւF�!�k.o�B"c˻�pXIY#�-�q��ۜY�^�N#z�AG𖜡T���$��M�R�8~�}|�2���1(V�9{h�ƍ	B=��L������M�yhQfn������W�Tr�/B|mV"��U}�Tkw�����8H��0��Ο�R�g����E]`xqpY�>'�%=W���c͎C�_��3%_&\i��*'\�8/m�^��j~<���/�XK��T�fS�:fd(y�p�$�٢RS#�˒��뗸ϻ$�,6=�=Wq�{n.���M�Jy9+B��'�Mh�"�}V�z�&��M��]�{�T�9ګO/��.�5��_^LGa��t�O%�&�$��f�r�Ѻ�<9���+]��|iP��_����'��ʥj@�����Ȳut��a3�}��ԟx�1*2��z���N�����yZ�s��R��#���Qu�����%
���v=������*��'GƸ������mS�l�9F�t��y�C��v��� �*�ْ��nM�Ko�]�e ���I�J�_I��Y��4L�������簲���*1.\��,E���
W"�T$���H��;���5�{E�}���ƙv��m����d+�(�<?�����{���!i�۬����gU�>_"T��y<�Ռk��B�ZzQj�Ϋ)�H��8�E�[r�����e{B�&ar�'Y9�Q3�j������m��剦4���n#qv�=W3�7	����[�ck�0�k*�|g��R�;ʙ�� ^f��V�ɪ�ۏ�����>���Wm.	�Q\�5#J��'���6�<м�ؒ�:N�%���K&N��\.��lr��sI9p�ly�L�.Ju��jѼ�L�yG� `݊�wf�١�����jQ�H��{�(�r1����Ӫ���V�&��N�>q$���/�{��`�����u�\ꌁ,�fY�;�wpa��p�I�7�[{%k��n�N�)6i��mV�D%sM��ðP�a��\���+�Nt��2`:��ӝ=tm�w��'�wXd���SheQ����l�+~�j|�G�%6�CכO���!q �$2���d��=_��Y�o�����8�NU҄3晵K�K/��O�x�z�r�4�j�F�q���B��@7�Y����B��=��^=�i������i�B�d��y��[�[ʗ�jv^�=��Q�90��G
!���d���-�MJ(4��*���c�L9˞̉�|����d����
G�����A�T����Ǌ!ց��o��<G�.g���wŬ�ٶ�;�6{��E�Nn��#yL�gg� !�����-�����EX�,�|�����K����ҵ�u��I��,��9�"��6�'�%��w�iJs�pz=n���<(��9���r6�ԕ�,�	�>��+8d���ŧ�ܬ�%�|��W���w��S����М�+Z�9���Kf�`���_��\�;ޗ3��u��K��\�Q\��p�~fZ�|���]g���@-H�/��x|��V?x�6ZC��3P��#��������zd�0?Ʈ�V��e���<�F$M�#�7�2sQ��/�B���)H�~�Ӎ�B�b����bT-��9�+�����ʱk4��F�n�#"��\/���x�e�s�v�)~������0)ߋ�Ֆ���m֛M�Q�ŸM��F��u�˧K>�����+��c@���AqJЛ��
�	ա�Rq>�� ��,�b�B� �}�����J]'�ϔ(<m\���_�)�
pg���X�;�s=%��[U���Tp@Q�w���Ti#r@�/d?�5�oo�l6L%�@� ��e ����.t�;�*avdȄ'��*�X�{���1���v��*C�	�W��y�u�����!�VV4ďx��������5\&Prs^s�x |�:��"~�zš�5����;�qx� ��2�J![.�].,t��}�-6�EV���MH��g�$鸶�W,2+������e�g���7g)�����}qg�2n��S<#�)�ȏ���s�F�[�A���Y�����3���v�� Q�A�v���L�mg�,���c"���;T��l�g����Կ��.b5���������žU�����&��q�����)kQR���q�wh=�յ���up}�8�w�h&n���r�"��Q'G��35�ryiَ�(ǔ����R�5�ߕ��/Q��������=��:���K�_)�6/���hsq�ҪT�뙘�./��N4�e�����ҡ/3E��^�`vP��q�gp1���P.�UH ��Z`� ��39���D�Iq���-.���YB]�j���Av�ՒՋ�����7Ca�L,���y��8�D�b��ղ�d��]N�
DNJ?O�_��Gہ���L�JF^>�qq
>z�I��,~��+��8G2Ϡry�R -�u�{ګ	kx���u��q��h��ocM���U[<�z'��L�滰�Ig>N�<��]��1��S+3����>S4�T�����*���v����۶� ȗZ�`�������ÚtQ�ɵ���͈�����M�F2����_b�=LD��2�E�9W�u� h$E�T���b�Sd$�}�)�R�4�)~9��)��w�s�l����Ņͧ�n�i�a��,C��_�s6U��s,�C=�骉��ml$Ʋ�(Q����Ӿ�<�
8��x%,voJ 0GdT��������q��aq0��K���M}z�o�����ެ�Ԉ�U�(��
�����'�	�� BUF�Y�<¯St	�\F� �TG@-��ռk���C�H�N���(&�~�C2�"@A���]6i����_�ML����+.`O�e�ӏ��#���Z$�k¦̬e�߱(J�������WF�������u_B�J<��g����q�V��ٚEݬ��h����#��s�:�n,O�я��ڥ��c�*g�U��ϙ_�[�����K����s�_��=}����I��G۟?��X�У��䨗L]�(��/į���uL�l7��I��X��'��?�I��7����=�2����	cKp��� �����׹l�Կ����O=��m�}N;�f�s$�i�ZN�����xZ����j���Z��W6f3����(7)�z�Qlgڷ���r��bNA��r�X�N"<�]�N��������5\Ak��J�ڈ��7�^z����L�$��`Ta7��&Ȗ��z��ev4|<�M��-PV�(zm�j�6O��#,��z:�tW�> �46|�V'����e�0���΋� ���s��?ߢGwsQ��Um��ܮB�G9OMCܗq�����%�.���&/H4���l�G��G�Yΰ\.2��Y4�?��Yҟ�a&>�:��jA��l��ܠ^�ߪÍr��t��R�3�"�s�+���(P�F�A?I�
t
,�g�xeX]� ���X�!LX��q�nB������GX�[J��xTT�q�/�l���/Ec.���A��Y�˜p��yuq�?�N��l��2�\9�^�T���4�vd�!&�o���p��h^Q`w����=�.�uJ���@��=jU)���&`��%�Z�|Ur�Z%�k0���9�*k#��ġ)�q��F��א��h�+�L�1b�6�F��ͤ�cp΋����=M8Xu$1���r����9;4�>�'e'gg4�dM+������7�][���{}�0J�(�ʎ�Y�����z�WO�S��w�G\n����4��Vzr���o!�����5&awd�d�s4��7H@j�>�P�;r>�6
�ؼ(k�^������X�~�bU���;0�m�P48�2�'9�ebGݩ������شD��h�	/�/����uxZ�'�BK��~�G����{�X:�
�jr�u�������j�����������I�Tn��9a{�22w�2=���֡0�^w�ջ��kӄ����E�ւ���6L{n=]�~<�eI���x�!�S�Nm�I��j�Rh�pk�6ۄ�rւ�����#㮆�r3�ܤ��l��������-S�I��"�F~E��۳�� 1�
��	T�bf�0�+�q�����|�Q��7�L��SO�Ll��t����N=ӽi��6AT`X��OGS����y�f���H�_�PV��F�ޱm����~?�Z*��uM��.J-�S�14��/
 ^�3�>@�Y�� k3Ʌ����n�CF����1o�\J�Q�4�%c!#���u�@{�S��̤�Ϭ�����El����Rtŋߊ]-�LW���w��Z|󻶝\���o�+�����h��m�{�%�r��]{8k�D�ѥ��D�n�(P��JA�U�|ƙ��RoF����~~�۷���݊������v�N��2���0� ��B�'W��r��Y챌=�G��ԙ�SL����I�q�w#��B��<c�'H�n�ai:j�����i������Y7+؂1���>֯F�`�B��9j�>�R�+�W������]��v��q��`n���1a6w%N��eӊ)3j���ܔ�)h��)K�%`���%i.l�{e= ����Z���Ѱ�D��?��[��Rjg=�O6Z�Z���"�4���|�i��3�m��� �]0����q�e�\$��P��ټzw����ſ��7ޅ�jǎ��.:�u��i�dh��	��B�>q���",�������~n�E�͗\��G�5�%�ɺ_%iE�ۘ�ƀ1H��m�%����X18;��G�Q��Ը��k
��֌�K.�ު�h����2h�S�o�����5�xR���(����F����cbs��O�e	�H��p��`,�4�/���b�q�
�g'�������U�e�:�V��\Ï�!+k�-�2�[>��a��z\~v�e0"z��ӻ�k�x��[�A	O?5I��Q*�|�3X`t�V���O��ŧ�d��Ȃ�r.�`�3[^��B{�U�Ӽ?�k��:�j�{�C0ϥd�@ o�)���G�Xd���^BǗz>���cas�9��|��H�:���]�������t@�W�gq-����<	��������Z��j�4'�ر��(o���n(����Wfl�T�;�_���/S����A�>��â* u� �^�^��ZT��0{�U=J��j��ݞ��,����z��St��C������}گ2�-9<��g�@��@jShK�kߒ��q3+�k
K�r�������t��c�TjN��k��6Lhf~�#R��(��0t��JS9p���8��d�n�g0�a\j����k�K�ωN�zx�=^�0<i���7��Ɉ�%7$��g��� #�n���<Jh�f�#����3C��Z�e��]oV�{���l�pA�hէk.�<y��oI��D��M@�������O�É�]'9��pC��~L_~]�a4�2~��=��$#b�M���R�վ������i$�x�~���Z9�Ğ!�^�a�R���Ery�ay��O��ٟ�����&X �O��%j��Q8���Sg:CdD�Yo�ps�E��vX@�þ�2B���d�係�)r�\�Kf!M�w�lqȓa;'��I��ti�(����s��ʦfj����A��M�u*_{�.|�U��`�Gd�N5*}{��	�ׂ`[W��J(*mSzY�p�i�})�{&�Kː���PT}
}��?�^���,J���¬.��E���O[�e�E��m�x�Q6��W�^Xh�UQ��蟝��r̅3���͎L/�Ki�8yvz���z�}M�?Z_�l��$3V�L��q��w�E�"������.���es��G�Z�26ٲ
�w��ԁS 0�1�����)�0�C�c�E�|�G���C����ԛI�ޣ���r�~���� �(o{	GޒmO*�s���-�t�P
�W'u�Y" I������vzPkE⸟9F�4�=�zl\`�n����o����vGKME���U�B��Q�s�Ø�nwu�]�GF��~B.1R��E�I]�ȏ�jz�CS��D$WvJX(�iRY�&ϩ¡���h��H�y&���Zn��*v^ʥ;f�);I�}e��vi���E�5*�Vʷ+\���_[���u�"N�-!�Y$콳���M��қům�IXF�}"}U���	GȊ
s��aO����OU��^�@���+c����xi��r�LdF�:�����2e�}��(�Ɣ�1��� �0?S�oӤ��C0l�\BC��w,H	�w޿��)k|�A��4�&;��b͟]�U���)�Ƅ_]! ���:��P�ө������	��ժ�|e�4�-���`}�|nXu�������e4��
u���?(*h�ʒ�n<�~،�������Y����JL���&�]���t��ȹp�-T��}�)��3�tF��m��b���񦨧a]&C�Y8)ѭ�)���ǧ+��"�v�v��WJ�V���hQ�L�4|s۩ie1l��'�����H!�u�_��-���Ŏ(���h�2Μ~Ȧ� o�����њ.�#N<g36�r��ۉ��1�朌Y/��) ���xbj��Ԩ?t��&.�Dta��d��-�S���B���|�a��J��RL�i�St�Af�o2Z�<��F(0y�ǰ�)�!f׫\��:�ڦ9���EJ���z&+���?wK��_����s�%T�r����r{�4�Z&:�����oY��f�#���C=��,�0A�zӔ�W�;�T��]c�b� ܈�V�Q�r< c���i6��UX"��뵟҉���m/��z����㸧��Z~��d7���R�G��s8"UZc�{�`-�w���L��e�m�ؼ�,<g������u�#�����V��~
w"L���1�ꂬ ;�����T��8�uz=q�J0�v���P*^Һ0�<A���{������<���7W�@6�}�bj�C0�I/�;x}��� Qd����{V5��6���w#d�`Ky��i��n ��t������4����>"��}�g��3��-Ek����|S�����(bC�fkcqHn�<Yp�U
�"�OZx��R�� ���h䅙 tD,�X���������U����A��:��4xO��@X��)?����}�/C�� �S��w���� �T��.j�P{�t�Uh_�Uw�0؁"�D�8Je�D:!���L����,X�m�(k� 1�D���D����'�`1m�|��YH�]Ng�Tr��jM7�t��/Q���4g>f#�w��CٙvJ�y`O�
h�6~Y�v?�����pÉ�솆�H��%Y���w,�>C�l�;(�aUg7(*�ZDU5��bP$��2�+�+�����*��~�*ufc!Q��<)@I��,r�nX�w�����\=��]$uJd�F��{'�Cl�he��Ϧ�����^ɧ�?�@e	��)�'�«a4�e�P�����j�*���q.��Q���C�Iv�6TV�. �p�1���*�Jխ��=ɨ?�'.n��iN[�0�f��n{BW���(RRĢ��1-ڼ��<UU��!�q
�4D����[���b���X#�j{L���T'G�^E�t���fF����&��/���xq��F�{��� 0�I���E�*;ȗ��ҳ_'n\WΛX�T����@@'��1����5�*�a\(��H0����@�J�\	X��sYTLE�YW�2H2؁��@�Vc�yz�=���fch_��Ɨ�o�r�F����fc����+���]���x�)�~��c�IFQXc$�̏*����Ԏ�R�;�	
"������T��U��,1�ղ��"ţ�� d��9Ș�z��;W��_숹�gS�#s5��0Pl�����/�������[�q���I�D9$����!�0M�H��V�8zg���/e�&���vuO����iY8.����G�d>L\4�▸���=	SM�^��wd�\���h�ٸU���e-0��K���΀�$E?H̐C$��C��K��5X��	~���p8�tW�&��m�SW2.���
g �)Ţ^ϕ�~���{(e��c�%��@" �m�������v"����ڒb@5�r�XS�n^<�O͚h�������\0Rˮ]w�`��JL��
߇����LN�AdK����s.5�B`ީV]a�~��*x�:���,�o4��v�w�	�+W�p�#<q��. �h�H6��5��������2�K��9��o������uǰ$�M�V�k���ұ��Rk�H��z���A��ǂÍ�	�;���AC['�̅l�6u�V��A�s�k@S���>���siq�6Ի�!5pD���`h��4� P+bNˉ���Zt���ߛ��wт���ho��`+<�
�����LG]5��U�|�R�X5��ջ�`����eO:�*d�[�6s\}d�D3�˸�U��\퐛:�c5	Й�Pz`b�hv�]��C����A��PS�;L��w��!��nq�@�d-zY�zԹ�V�M)?��Uy\��G��>p{�5��ɼ�U����daed$v���q����:>��F�"�1�\��f�.�y�����'�� !��gK��֒eynm����aBI��ު��v�n�d[<�&��k������#���^�/R��+���!@w@�(�B���ݗߊ�Z�ݯN b�����ݠlo/ɥ��'YC����*D;����茙�:�VUQ�ž�f{�ߗ��ނ�@ ������ߟ��^��7����qn\����+A(�;TjS�p���@�L�4
�W��/G����!�� (���if�/�V��t���+�Ii��|�`����
�Y�y ����RΕ��������@wx�Fc{(��\F�����'8Չֿ��Q�X��Qp�j��Ef uHkN�m�e��]v�"D������4����h��[�e��r`��7�����^1F�kI�	��C��9�s�m��Z��Rb�"N�|��_����i��A}*�y�����ж���6P�Q� �n\Z�7H����5�1�{L?G�h���|p
6āQ{r��s������\���d�!3֦�'����xc����Y(QX�\g� �J-P����ץ����wc��]�(�O�}dg���\N��֏-�5�Ko�"��*D�݀����Lѷ�<��w@�8���`;+�۸�x�F���n%����o�q$��9;	�§���G
�c�."��hǊ��6�%��>�D���Uh f�`�v��������`R�[�;��Oh}mڒP%>v"�2[���N5C�'���HjE�o;��]b�,	Q��k�����J������v׵�ǀ-��_V�2��M��=澉�޾�b	���
�>���D2�U<���1�
����B��L�dr�,΂ȡq����WkJ�:O�gC�&f*�L�e����<�a�Y֦���h��Z���$��}�y|������m�ȁeiĂ���Ojn�{�jA���~R�֛e08�!�({���.WLB.�mx�U�
 �� �ҿ�Δ{�H����Տ����xc��P�8����5���j�V����"��OV|}��d� w%�>#�]�����=1bV���h'_�=��ʫ�4e���߈��b��סGgأt�&tk��ֻ�n�QzG���%s:)|[9��<�mu�-����gA��{�h3Z*��z���,�[���!�,w8բ\�I��~R�B)��!@��אPU����^�vc��+����(�:����.� %��hQ�3W�/�Z�,�h1{;R�m ؍��n	�!���o&�t�4,,�7�A�1{�+���%��R��$)0�5��֏<M��9^!*��d�����WppM���4?E�� �7Sy������U�1�q��N��$�����u�N]'����1�HqV��>J7I�TI��^?`;̮�J�⛠���N��W��2�"�I�Tmŋ�y}1��1K����V� �\�ɂ4,T��(]�`,��u����״��L�4V�S�++cY �>ܤ|�nVg�/�y���Vy���FE���?pq��V|$�}l7�L�g�{�����+��@T<�����Z�����ؓ�����j�:f�9I�*�z���KV[�;j�{�_�?�"�9qv�a�O�1������Xr�^�s;�H=#2�c� ��ӟ� ��r�0>Q��������=��H"&��~*m*,K1�
ٙi���K��YU�S�1,]���l3�x�Sp��������?��=���U~?*�'rQ��}6l�T���~�P¥9�Wsso�W�$�Jj�W'FC�Ϗ[���m��&����p%�^V6���Tى=��M�`W�ܗ�2P׼� խ<\4�<{���F���J�i:�I�	� aG$�e>#���-p�EBp6M�K�6E�H�<�l���i�]��yt� ������z�t����]�"���"R��	�����b�u�@�~K�
 �<渮�,��R����5����sٴ�K��d��d���vc���@����)���z"����xZ����t����~!�����?A:UR��-,n��ׂ&�.Aj����c�܇�zl��v#B��3J��Y��-�������ְ}��`�8��z���k�Z��E
)��R�ׂ�Y��+�
��3�0��N�*�?��W�Ҫ�Ď��֕�U�+��4���s�:�E�:_�/y2�����)��i��`�����MPx���E���g��d��JB��Kk����l��.h��'\0�ٝ�}p!?��3�Tȗa(�wq �F�ht��mm�V�r$����JV���Z��v}��f#�П�n�z.Q�9�"&j��+�.�F����������� �:`b7b?!���� �)�>���M`�L�I��<�;�����1g9%L�1sn.�Ms?��jM&5�a<�8I�nm��Y-M�S������)o\���?��^��e�ұ�ac~��lŭ*I)�F5�on�D�#��i�&j��@�9��ԭ3�w�Yv�{gT�r��xG|����>��T͹��
�����Q�%u�5u�t�YJ���1 t������B���N8�.��G�O�.�A��Fߘj�n'���&�5�T�E��+���~�b�9c�j��m�@�wr� ��?��=�Ls>�Tic���ӎ�=t�c���A^S�(F�?�J �~�Jw�����&�Պs�@�.>?N'���*S`�gGQL%��s��TjGb�A�ǧX-顄�>��5f�؂C�V�Q+�	Q��qyT�u����54�Lu��[~�~
�_��wG��w��`����;"��SDϬ��!�>3����m�>94�1���R�.��S�U���b���vS
�7vث_�fdO������gR'DJ�Jl]�[�A2���	:*����g4��o���P��+����)��m�}{��5�>6Ky�z4s�T\���0g�#��#Ix�<�|JJ�>,�rj^�]�.�hyw1�����.]�����.�L�%|+����f�h3"R�+��]��#��O�hiǷ��mܻ���u{��6���k�У���3z	�i��nJ��H^�:�P�>��8�
���R�)8��z�z���<a��j�%J��|��.�I���c��ǯ _�M�c�&jL���Y3M@(��P�г1L?�`�c�h���)��M׋n��g���Z����9���Y����-�+`yX���QWx#̜0�ִPC�R:��k��.F�GzlQ�^w�K��ì��;c�*̯����e�u|x4mK��|85ٚ=3���W9_�uL}W.��wo���>_�I)��k'K�2��Li���a�w�1�������;;u�w*[���E��@M��]���Mj��X��zW<����p��`k���-�~j�����Mg��H��mqd�+��y�����j�p�
).vc+Q����N}��-E���q��џ�G����,�K���n��VTH;�G#�F����љ�,���;-�q���X�I�3�Z`i*��V�����RK~�JT���j_�VFG2F>h��6j[C��N�=s� f�J��:n���FZN"�6�rJ������PS[�Э*�/��_�Nw0�0,b;�����o+�Ȓf������VY�W�v\y�:J�꒓ƃ���NV?)`��RaI�sܵ�.d�fz�w'�u�^�����I�ߤ
OZ�����]+gyD���i5��0ҐX���>���� H�~PlTN�s�˅ԩ��I}�L��r��}w0%p�;�ۍo3�4�u����#ML�hPb9Y������-��#�	��� ���P6vw2��� �yW��'�d6��m����.}����5-��C S8�����;�xF�J�Y6wnj�G��Yu�y��U;N�\ 8��C��"��LR.D�L�)��޹/���9����0K��[��nE
��Y�~p:��輒��f��q3��u��E(������߷E��V>;Ƒ�Q�w�����zRW�n�PZ$m�:5/J{*?U8j��),>>�4���ޝI�
r���a)������A�q�)V�^�M�y#��i��lp鰇��/�^��`@vF&��o� ������~��,Mo,p��~���@��ae���K�8:��`)��G��&0��:�/��:v5d���G��ۂ��zm������K��X
��R�>�,hiD�ca���ӗ�ަ��I@������/�/KW��i�yL��#O4�W��x�r���0�oU���4Xl��D�.�  �S�Bmt�_�;��a�@�C9h�~7<}�*�P�!�u�ǭ�<����$��K�E����A�m9���P=��L.ɀ��t�8�Gb�#�N,u�yk��`�&!��mTT1ٗВ�*��[ �y�ܹ�k�cJf&#o/�f�a�c�|�i�$�XȠT�˭����J�R����ܘ r^����&I���H4̻+�7�OL�������"[��_��`�l�}�eh��aY�p����Փ5t��D�?$�<yQp�OH�E�@=��@`ħ� �=�E>7��fI��J��?h�L�Z���
G�
(J8>l<Ai{��zW/Y�'~l�W���0;�W�Ej��r1�WE���|'�d���G�ӼW�<����u�<�6X����	�
�Z���Њ�?���	��G��_nCH�DX�����g�B �$�^��B����zB_�-�-7V����k2�+p�'sw�>�?�:ew�+b�% j�(R1uEd��e�6/0�\�P�f���=�征�ER	E[
A�v�
��<�I+V���W��8�hK�Z���sO~X��Cts�#�~�M6)�E�&���6,\K_G�%%u��.�n�ڋ��{�
˾o���&a�VO�����1��2�ñ�{e��;���#X.^�7�����M���o���:C,�m�.o��A�&{���gl�0�FQ��E%��1�)E�rz3ߖn�	'L�]�Z�,�����SZ�x���k�	TL���!��Xs��W��ߎ��ߤ��!��+n��|IX �q"Ǌ��͑:r(X�h<V����>���m�Zou��S/�h,��J�]��#��~��R $2F���#�HJ��g�"o��/T��&�	��uB���g5QQލџn6i���,�^�7f��֎����M����zA-l�if���`N�d�����%�2tAT	� �\:!<�8���fq��F���F��,{�Fj�'R�T~j&q�]d�N.�@T"#�n�6�3�P�XĩS��<f3*|��^��O ��zx�$�(�o[��*��9z2�r�;}!E$wŞ6�L�Qׄ����o����PZ+3}B�Ynd2��0p��a�,E�m	Po}^s���{uF�\�v����
��/'h���#�j�r��=|3Gˑ:���0U�w�� �R�zwy�<�X��B���%IF�>&z�9�Ipا<������̕��Z!O�pfH���?�9�5�Ѿ��VdG 3.�/�?����:��I[=�O5/�<�_�oL\�}� ��`�����Aȗ:�Nv``rZ̟#SL���ra��bKPb�td�쏂!_�F��g�q���[;�S��ʕ�#ˡ�t��B�dv"�6f��<'@�y�T^~�Y.�>�R]����},�z6j#b1�'�g���jm#�j��D��Dˉ�-�> �=.e]��^.xys��&e׏  h'��S�y�X[!�����h�������d�����l��'M>�qx�~�����"r�lա�����%��^�ea�#�.���y
|et�ƞu�;$ Z;@nƍ�	aê��r"K#M*)��K�N�p���M^�KN�\��*ks�퐟���'
�ߦ�xO�RO����ˬ��w��H�X��\ͅ)�`�A�t*�Jr�8�dʍ��s���Z#�+�JW��ެ9��C�d�Y���
	��OJ	��3j,wD��w�zW��j-E��8P�/Y��w��P�Ah�7��<�1�~G:K��{/í"�஧8��L~�����sE���W9��f�@m�"�r5@w�l�:~v���2O����m��KoE$��"�-#d&�N�%Z�DIk;ܘ�.�-(f�:�ܔ�ϲ�p�}V'༿_�����D���9�g[�3�mf�ui���eK�.���$�>x�C>`�2��r��:I��?]tP���T�e�ܲ�=�_LĬ����?� �P��v�� ��yd�rj##��*�=�`��F���g]ˎƌ���Vg"����|n��A���!�L�ೂ*�`�ZBة�[��e�'oẃ{��Kn�j.sΡ�Ry�m�/����柗\ب���\�A����xX�ɐ��r�	�*�I��i'��7;z��C����i���{?�&��>���xB(�������L���"f�]�⚢���8�AtO�����	B�H�2��.ӭ
��E�P,�v��H��'L��9�B��M�Ln(y��`m��(�>9Ld �0>����ق,��࢏�
:O�xK�喻�#,Ve����� �J&�T�ٺ���v���rP`߹���P��*��5�TCCr���בyL��W�`��E)��B����Px�)��E]�)#��c[�gk�D;G�AL��N:��g��T��}`�*M�iӜu$�j�,�\^������]�wk\���^�U1
�vh	�8r'r�ɖ}�6l|I�Y��,l�I�r��a0�����_.�څ+5����e���2+�V��S���߄^��9,�K�4\��n���(])&m]콉�l"��������ՀR�1�M7�&F����&�[H/r��nʻ�%~���-��G[bJm�z����U��i�K��ҡB��6�X��&O�W���qڤ����hl�:p��4�v��[/�5�
q3XOu9�#@��&r�+%~j�Ӹ�<��$d%%1A�,�5�Z��Qn��S.^���x�"}E��x�[���}�k>�o5�L�ٯyOO�U��-���
�T������d�������s�!W:i��	�07vp�<�_C�]0*��:7�ׅ�`g��C����b[�oO�g{)q��Z>�����
��v<�̘��G
���i�����6[�`(E��V˖�
��Z6�MW^KI�jʴ)�L�;d�њn+o�0�mǶ9�ש�T4+vt��nc���m��ڹS��!Z�@����(��j���x�!d��N��/�;  )��T��z,� ˢt�	#����쎔�A�_5� -��"��S�ԩ �mFysdZ`��p�B%�h��Y��%�^Qg���kq� �D3��7�M��k��P���\Qzn�;���4�L/őE.��7�m��Kvӯ�7��,�fACe�|H���2�ssV��|!�v"Q?).{Ί8����%4�cg�0��	�ۢ=u�aNw�	?�:�Y�J��_�@>)�����H�.�K쯕�NK��:��v���%̚.^pʗ/jko�\}�@¹n�I�./�|>_"�j��[.B�������<.�N�r ��#2*3[)��ob:�!\=�ݼ���D3�Yf���Ѩj�?槊c�lY��|�^^A�b��/�x�y�����y�����܈��+�56��W@qG�R��NJYm�����u�R��cs�����y�Fw�H��OÃJ��k��J�a)�dp��}�X��?���as3���xl�IQضmU�_��l�4�'j�o�IW#�;�x*(��r��)#�,���W���tq_i=�=���]���ң`ފ�oF��(t�q�J�<D� ti�i𕿲�Ks,_�ܡ�W���
�Xح��o(Cjzp6v�/:2*,~��ѱo4=�����GOc��fVwD���ut�/R��F>X���!|;��̗���71�A���]��L�f?�@�/�7��Ĝ����t���振PQ"i��$�]���K���1�bb)R2�G\����1�Eb����͔T�~B>�mu,�6�vL�
�80;h���W߮��Z�̣�{H�(��ր-KdZf�2Q�\�SL���/��R8W�#V�w�1AfD}�L�,��mu��(���
³6x-,Pn�4�����>���w0���R�HK�\�s�u��[.�:�	��Q7����&u���X�Lrz�Gԥ*}ٷ�K�Zm�"�1��������;ωC���
�P���I&J=����/��$ �hZLz��"+�q���S	��y\�����Z�6$��J���@�4WO8�'�d�`<�`2��c:T�(�*Yc=ݶ�8z��-"��2�{��ג�4m�"z( �].Q������=��g1�E|f�6I�i��Z��^��y傽�),����XY��}��d
	q!�n�,��b�:�Q�y�8�7��;�0��F�c��U���1{�&o]�,{���q}�G�ڧ��bsM+k���)Q���4�-['�@�UȏdO8Q�.M8�Fc\��K��9��y�����v�Q7A���(���n2��$_/!-�V��B��~^�%&w�z�Ac��%� �ʡ��̿�Cw��!O�"/?T��Q@<@��@,Ł�R뎿g1@�B[O�J �Ίt\6ʿB�zꅌ4�,���<GZ�Bemܧ\L���	����ʂG=5n�En��m��J�7}�.6���<� �z`B�穧gMO�LKWɢC��M�����9�LXW��*�"���в��wo�O��2m�C��3���,�ژA�3p��s�8��F�CKwI��[J�����-  ���������RN��@�	MAWrV%įa����EW�T(�_)<~����������N>������r _|�`u��o;�E���d	������@{\Aӝ<���qWdc�����R;���"P% ����f���ϓ���k��"];;fg'|�Hڅ(����,�h8Q�+��蝴��IԳ7{X�S��Jv��&����T�Y��G	c|��r8�Rcx��28~��$�U��Wv�YV��T����HCL}N�`�W��H�+�o�NX� ifPu���l��Ÿ"`@Iy�c����*<���2�*������{.�B��-��^��:�٤x��/��ۡ�S~�N>��ˢ� �Z��7�Tg���ܾR�*���=�9��[r������zVP�����b�Cʉ�Ń%�ӿ��d�+�˱�	B�U����n[�c�Q�(X�o�$s?X���P��L������%���� ������J���6���l�/Ì�Ž!DHjZ��R*�z���vk��҈6��<��`���cN�=���(�//,�U*=�Aw����0��pRK���C��0A���ES?�6�����e�ߵd�s��@�AK�h����ކ�
g�������(��%Z��u����#/���@w�<�R:j���<�0��������)nD�]Qǡg��޼�͊�Z\�uT�n ��H��B���V��[Y�g����x���:.H L�Pp]�h�{	}���h�S�~�͕JP��dƍ�O�!�9G��P��dZ\�~|S�-oܗĪ$,��5�J�C��Eae�X_d]#i}6�Էz��U�RKqs��@��*�j�+�'	�U���*�U��Ɇ��%D�\��[jZͮE"aX�[�-꾛 �Ίf��6Y��>�FI,��<��q��Y�~s�����Neƍ�E�T���/��KZ� W]�䨲p`oN�d,A�wt҂8�w^��հ�N'7e�)��I�ˠ8�a]iζ�D�Y�������[�n�[��͟�}
�>��	�%�S�-��z3�OAH5!6}b�\G������04�4d���������V�,D�����kZ!�d�i��4�풯�w��io�I���Z;�P�g�;4�y����0W��Y����1t����	����E/d�@���;p.p���|A*qU�oN����f׌b���+z�aD�Q1{�>pP�Q0ΰ?��Um](�_^~KihZQų��_(�]38�i� �;�4�Ԕ�ĉd�6�j}�ܶj|=��!u�B�Ov(�n }������>���E�T�Z���`@ִ$�!�uߐP 5�9�1�u�%��ǚ��_����#mt�`U]�IR�K��>AفEl�r Ť��h]�a��2jPп>|l��.�OM�Lo@Ig��g��P�Ř���yR�c��r�&ؒ�����Z����{1�Ā?�d�UIH��l�zW��Z��Gʇ_����"W$�ʠ��l*�C��zT&�@�ulﾀ0an��Z���Ψ��Q�]�G+"'���8^N�hJ�.:��#�{��u���wl�L���EKݰ�t�tO��{fɴ����j�x)?�h�sb����X^ϙ6�E{4o=���"��L�ÿ�ix3"���O�R�v�����(�X+2P�g-�t�Ө=�\b��������cj�͊�oѡ��Q����M�D�7���1�?���5j(���_�8-]����l\��h�؝����}ՓE!��jK	��}�F���*w��yLd��Ϸ�Ʈ�`t真C���k�2�x�A�겊	N:0�W��Z�F���J��-�_�X���i�pAG�`�Ǯ�c^C�F���j�e_�?�ls�U��Ż=������-i����f���2y�x�d��/kZ�+:��+��w�وòaB>��x,�v�T&��Z��8��Ӱ�Q�E/��t�Ϊ��d\�e�>͒Qי�5w�E9���ʡ�$w0Ql�&1"[� xj- c���$�i�#`��>���bԶ��Ө)v�rۣ�v���"�'1�՘�9�d�J�d֥�+��@-��7�{�$ip��<��������?z��<Jf���g�w߳=,p8�>�rdI�¤t
d(S�-;���o�d��B� ����bW$����b����� J�^�QHX'� �μ�U��kf�:���=���UO�l$V�������B���[ڢ�mN�������Y�:K��/����FΆ�\�*����E���!�`!��ט\c��߂�fem���,��ª4&�⢗�E���%��?�;/v����!�1Z�,/�v����*v�xq'�5���mfZSJ��`�.Jp{R�E33k���B*�D籷����lyF1���Ȁ����'�Iex���ea�1X�Sz�������ͅxy��G	�<� �1(���Ɠ�R@ �,e1�9ϲ`�^��������~�
&{r~D��)���[ ΃K���e����W!��H��d�b���'5�O�b�M�6�8v��SX�$-�u�&C��s�E p�j�k��x���c5T5����`>�Ý�Y�w���m2~���QeKK{m�@!x�������]؝Ɗx]����D�җ���1t�aA��ԧY�F�n���4`7�o�����Bч��w�A��l0���q���.a$-}Mw#_�s����]Q��A㲄%_����<,LǨ,�X�7o���u�d�P�*W���Ye8u�Z�$���e��j�K�9�
<���G��J?Q��Tfpb�&�|�L���xW��7m��;&r����w�����-�o��x��$e��~�ME631���n(P.bOd<�5�J�pv���$7ML9�zih�3����Ǧ��Gb����� ��n�h���ڋV5j1ӗ|����l�S���9q0pϣp�m)~wm+?�Y�!�*��0)�R㕻�q[X���{��6�a��E�ʥ��/�Ⱥ�@���J����u�m�{�����X� �<�d���7bs��.��(LK&�:&��r�>���11���i-����؀���Щ%�8vcD�mR5l�v�ه�;p��/���'J�OK����昧�D�� ] ���O���cì����J�ؓ/��#*ş��x�W�:Vf��M.���������)^�5�A��.���1 z���K!����Oڌs�r�����Jz��b3tn����WW�e�n9�����ʥ�9�d<p�� ��18�����QƏY�����k~�#/PW��ۿ��-��ħHwɲ��ct9�G�u�]d��x!+��Gn�Љ�7gNӏ4݊��L�3Nqd���q�\���� rFv����:_�ƲxKf�f~��[��G.�;�^wL/ l�ء�h`�c���-a#��}Ā-#�̗�mj6Q<��kQ��oR����q̌}���sA��)M� |=�$/��-~|��b_{�=�Q�e�/Q����������G�P��-g�@�M��۬<���;��jzҳL�$���rc�h\lX��R�k��`8����Fs����g=tu{w?�7Q���n�E_-@��"��L6w$��^�50��B�߷�F�k!%���w�4�ŞQ�-��C�>�N����O�K��8�I�>ݢl��D�ձ$$���̋>�r΍�'�.m�2����	���ߜTģY�mQ�?�zM�*-�!m�[�q��HE�~Or����D��3w�-���;��Å����gE'1EH�jz&�ܳ�������X�������D�3m���J��o|I\B3�.��}��q�[׆�(�0�$�/�N�zQ���ꨨ��UdG<��K�.�@�T}s�;���0��Nc�E�B��ta0��
��	d�1E��U�[�b�E���k�E��� �Q���Z��jnN�f�:�f�*�� F��ŉWAt�3�U`�ϐ�v���rYǜ��/�J~4Xd�d���/@ `��魐��M�lOwd������u��?��bpg��j�`|_'�[��(��"Q�@O���
<Ă10v� %]����W.�=���62�i���-e�W�E��ѥ�v�w�Q��fd?x #?V� �@0���;�*M³��r&-���Ɲhq~Q=e%'��D������˛V�:Rt
�5�J�"�L/n�/�)���V�$H��@$ҝ�Dk���$��2��#[(MHL���20;+zQ@��B/-��D�2� �s��p��m��B�2��Bi������ڳ�}�)MAܔ���l٥�:��T�M�e��␱(�zߞ�껐�����W�A1���D��� %�ޕ�X������C�G!c��������&�=/8��������8q�!U���RxM��>	�D%�j���A���nڪ�[
�f�+�es����;��A�Le���\��fg����$m���_�HKr}{0��ЏA»��3YwI8�����E�w�>�Ū�8X��a��|��*�Eʮ���	�H]��ܿ�z����u|7S#��e�`k�M�Ym�p��쎀�$G�S�)��vGDE�<B;����T��[GR�^��xK�M�+�t�]�hJ�*�����}m��܄�'0�p�"4u�ܐ�=+jn�� Q�fҔ�x)�	e� h���=ֆ�_��~cX8�_g���3?�{u�3��Ό;2��镎�M#wS�+4�����N�cO���@��)�D�?E^\�F穕�Vf������;�i�`30���a"�)��Ś`�U�,3��+��������<��]1l��n<���MV���E�L�^�1O��6<P����P<x��m��I���<�I�%�9Rw����H�/�m���շ�Q����m;��Q1���{� ��W�0��q��S��:�R?$C�p�C��F�:���q��7)@�
�5¥�-����ҋ��գg��w	�X��h��k���4��S7/������P������[?*s��G��Y��\۴��0��H�b�R�2|	������Ӂ	@�H�>�R:��-�kK�B�[j�5�ѝzy?����a�-�+����f��+���&��YBW��U?� '��@��/;��ҼE��p����\��X���L1�G���Nf5�`-C]����8ەw�%J��f�!��(�\v�c���o|��$��h�ڜV˪kr��<ĉ;1?u� �ă��n�֗x�S$AL�SNW�!�j��`�<6|�*�����S
�w��N]td�\+���.�h��~���CW�/��s�R���d"9�K/p���l�w�n〆o�Y�%�j|s��U��*�ʛ%��AdV�GBC50sh��[i?;��� 7O�MrK���3���K���Q=2D���+�ֈ2��i�6��YRRD�Z�Bg�YJc{Lt5������p&l��9�=�>־�R�V�p0�مyG@�œ;�~�s��j=N*��U�IkG�Im�U���ɎF��`� %n�5�]��Ю�b�j�{e�<>a��o�/џ}��b^���μ^l�5��hȤ�8� ��i)z�����+�6e�@O�O0���x��7X�V�r�Z���yl�a(^��[��J��;�c�^8���}��.c׹v��~�=:� �H�Q"�^�G�8nM��*�G��db���{�
�P�������i�T�v���%�o��r��|Q�ܫBS�P�k���f� {��\�o����ڼ�� ���Ͳ�r6���םiJ�ͼB?KF*����-Y%�Sx89�{�t���G�'$�-�Ƃ�,qo��'ǥ'�K��U�	�`H�� �X�TR ��!��R	�Nb�}�������ĵ���	���P�y��B������@�ިpG<�.��8����r6��\�p!S��u�P+'3L��~ByE��jۦ��<zt�ǚ�A��w��"MH�;���LC�Z�K+;����H+r�d&mR�����K��0a�X�2-��KD�Z1��ۼ���2�7 "���**�Ak�mSS϶�1W�;�1�־�O�yW����N�m)L��
Go�w��~7^i�w~�;hDO*?$��,"ޫdU�\k�Y7lIKESu�Dw���Ȭm�T�,/�{P6q`�+�1��D��C���9�6�����n�'Vo��;5t�RaЊ%�L��
M*@���]�킧�� =<�J!μ�%C��iy��64��<��P�}����0`�Q ya������g2ƣw�J5�ߐlog����uDY�Wr�1̇D��0Ht7��w�P��V�M�$�e���]ډ��h\xN6m*s!����g���P�%2l"I�F�e^��E|ٷ�L,\/yXS��hX|�1�[)�Թ+rk�'�u�u[_0:&X�Lf�S]:�v�ת	 ¡ܰ��k�:Aʝz�fRo~k��7� ���Q����;��������Z�@�>K���0�+��W�D�_�1^fm�<���	��5bMg7[�×��ێ2�p}c��6���F�����--����'�ӎ��L�@
<%p�E�H�j2Z���7�½N4�-^�~ĆoBG�))Q�Qk��帚e�e��5#�֏��g�u�O�fV�  ]7Jw���s�kĻD1���a��)l�U%�#h��C\Q�c%�%pa
��m���Z^��U���Ȗ���=7�q����NɈ5���ij�O�!^/d!�Y
��Db����4]�X��mf�r�����+��׃ڜ��!	�_>�V"Y�(r��$(�u�0���+OgtŅ�9�^UZ��DM�˨����[ *�!W��K%���������ȟ�؄W���ta�_�HS�'t�(A�1N�Rȳ�?ՏW�Ro�� wGdba�Z��d�O���beD�6�"�� �.�q�91��*�uwڰ+��O����w��fLU*�*��ñ�����dT�Q�i���TH�7)5�Z���Օ���'�5z
h�VE��C:^�Y�{k��s'7L��A�-��b̙e�4��Hw�>�&6�X]I�a�/){�����E9q��U�<�bTt6�ĸ0��?'��Y�/'&��1���F�S�)[!���Ҿr� �:7�f����^����(q��<j��>�DK�r������'�V|Pq�����q��O�	��t(*'��yĆ�|��V+Vo�����p�o�����Xh�#��|KZ6�H3go&6��'�.�KZ��;�0VcW�z�<Ϟ	��G ���"0FѼ5��$���(B\ޛ؂�|�؛׵���7�m��Ջ4g�%a��H^��s&4<��H���VR����_'2��֕ґ��s�gɟN�LZ�<_M	����k��#�v��ŧ[��U�k|����a`��ԯ&X$��T�[��@���Sͨ����w0���{ ��*�0:�����j_C�+h$!<KɫJn�;f�p�6�wa8p�](/���u�NG�0�{��Jق!���;'�6Xg �E(����� ��)DK�$z�����P�"{�T� z�6�J��wy#L�ȫ�!r<iy�i�kW���s0Ne�b��#};����`�V#�\�2��?)�J�p��C���;A��1���v!�>aAy��I'��aV�&��5GQ�Iy�M�u#����R�Jb܌�T�o����3�Q��&XO!��7�-�Y��ؔ�>S���1�hv���u�enm�����
Z	B�j�Q<d�`>��O`�w1��@J��L�?��h��±�}$6�9ȴ淖�)�v򚳪����G\��}C+����y�GrE��EUPK�]�����Quf{0�6�ّթn4�%�̳_71�QNT��@�F� )
���/3��+w��ψ߆�y:h�0yw~����"jwd���#{q�1a�8Z9��h�> *�ݷE�$�&4l���0�r�����\ʁ� �.Q�����#����w��$���<���ҏ��Q%��J��s����z�YB�[t���Ł��otD�4���%��1(�\���fT�$�y�*��C�,�IkmD����n�4��k���T-�"�}�L�|�����/���ԑ@вtr �5ے�W�����޸ʾ�DV)�J6�s��l4�{zP�zÇ�_=Z�±���m�RDN�(��Q=*��&�|���M�
E.[�Y{���������Ї*(F�]��A���H�{�jD{���H&.�/mz!�<i��(=̷U�m^���#��chT8�`���FhR�:r�H���K�g'���L+@�]����*�� ��=7�cz��ǩ7�.O�����J"��xR����J�+�
���f�1�=V�]��aȭ]��FS^[]NR���qf���^�����Z��^�i���i{/�<R����-���˟Br"1^�לF�.�kjz<ܿ�E̻�C��"�� w��F�XH8�ŢBM�s�N�����]NPr����p�,b�'�%A%����Vp`��`y�!�Fjz���}7�*I%"ϟ�@��v�PI>
�T���z���bS�QK���2�F�&H3�P�h,1V��&]�����i*]��	���!'D��x��c���%b��f 	"����<8	�04;�|�I5Y� |�P��C4�<%��~+ؿ39��И-�t��s�v�2_�ޤmQ�z�E�=q��F��YQ��TI{�C<�-�S���.�	�gl��D ?��By�Ք��x'W�~��mܬc�;r�:UEh���v��V�����D4%��:�V���⛔��8(�#�;��K�<��@�%���0�^�u�;FS7i����A:��X��<�O��D��*��`,�̸�Z�?؀:i͡��Mx[�4���|訠��\pnk����π%r���8;jp�~���3���{��5YNa��6hza|Z��C�'���]�D6q�a�/Y=�y@�:��v\/R�0���{�f�V��<��)�DV��@-b�-����R�qI���VB	I�iU[|U�-)H�x1:��v�^Q���-�H��rbn\�ސs�z8��z�������$x7H���k�	�h�%�����5��3�|�s�[��<�͇*:ؤ�?.���*��Xø�7Dȯ[�c��$��/��4E��lC��a ���g!��;��Ϛ�^��R��Z��y��v���j�CF�	ϋl$	$F@9pe7��u/�%�ަ&N�\�����N�s���\C"mK[8T�!��z ���Y1E��9=J_���Y����İ�&� �{�ڟ[8�nA�|J�7�W���W�4z+l���$�(D�m��3�����y<�0����9�蓚��O[Ԍk��TSf��aZaC��O����t~����2�1f����G�ͲT�T���nh����*�}۟�v��G:D���0�lO�S l�Tw�pp�Qßy�Q�ˏYg�aq�r���	:s����-���ɨH��[d9��na�����\F���:���*��[��T���ϣ����C�4��	Y�)��jU����l�ت���]6=��'���]�\�|c����4vN�6��!2�LK�����mv�r�I�jI(��4h��F�uv'}�Z��Yٔ�ԭr�Ƽ9M�|��}�W,TJ�m�!(9��"yl��{��r��ةAu�ģ�/� ��>�h���cԫ��}�'��Б��U�}|�<P
)U-��w�O�L�l���`b:|�H�h���Ɯ�S"{�zn�H��
yv�&�/�oj1p��&l��\��aH�-\����ֳFD�v\(��ATF���'5�h"�E�H��I2l�S|I�rI8�A���X��>��:����U ���w/x\���߆ڋ��R�kG~�����|Lbcʬع_�tb5�xQ?���T"d�+�E31I��bP���/9R�T�"�����8L�Nxؖ��Z��6��Y��>���Qv����7��if��;H���z*���b��p��O0��A{$��`C��4���L��V���.Փ��1,ȳ���lFD���������g�G�;�QX�'��pJ!1��tQX[�{�	�A��wO�)���_�ܒ�I�Tj������P0��g*JV>:r����Ǡw_H��35(�M�QT`�܎���~��$:6�X}��J��U�d��b�MNN:��p�����h(�3�<������*	��_&vʡSƌ�E7�6���Q��f sK���� �++w7\�t;��������a�=�i����uz�U���'/�^bJu]\��o ��=��/
��]B�;��\&��Z
c�{"Q[����X'��P�I��Rjl���i2=`����Zhی���U�$������d�<l�?�j3M�Rc��n��#�����6��tlq�4��<�rUe�!2%�'�Dr ?jhG�<M/�>~��]�5ne���m����7Z=�#`�"�p�v����;�F�@��t�9������+�3�zW�a2ΐ��o�����G����,�9�<{��ʢ�T������c�EB�a�b�ec�p���Z�%&gX̙KG~q�H�xzʖ3<��ʶ��5*�0��2�9��EK�!Ž��l��R=�(ѷ�C¡x�6���R���i��2����!�oҿm����
h~w�R�!�G���,�'�$o�
֖�=��q��`���Ӕ7�c��b�`r��h��we}z�-~�I�$�tt�Z]����$b6Rc044:��b�{B�?�ֳ��:+gP�H�����[F�P:#@)�����#���;���IJ���2|���Z�#�D��J���z;�{�
 ���)D)�����og��1@6�4�
s��1;��"U5�x�9X`�pa�b��;�Bm�\^h+
^���h[�a���7�/UL�߷�;���w#`����?J�p��Df��������k��Q�w�����2 ڴo9�:[���<<~�J�/cjp9{�b��>�`LB  O*Ml�!�=���(��qW;h�)>R����Q3���cy=4g��oQ�pR �	���WV=P��XG����*�ż���Si��`���ժR:���8�#Z��=�ԥ�y���Cή
�hl�S����EJm|��SD�mZоP�b_�1n�]�'�Oj[�Ȫ���͠��\s�d�����n��d���R���!B�=j�W��3�jϽ�ծAV�Kӛ_��*&*Ң�%D��?JYs�JQ~ ��~:A���<��C�s�%WH��BA���lXh�NP���q�
]���Rg�"�uV2��ނP��7�i	����̵�8=�U/e�۳��ָ�N#��~�2%4������dXv.�e�E���3��`����?�Ȍ��+O���蜵�;'Rً�'��F;L�2�n �PJW�m	����q��G��� r��;�P �V�Klǆ���{Ő���&*�*Ƶ4��ⶶA}`C2n�}��1�Tɓa���!;v�-*J$��j!8Yd"�6��$!�8P��85��J	���V�̄?��D�Ԑb+$���÷{h�r�m�9
d�#���{{5R饆`{��#���̤���$#��|�����S���Y�H������L)�Y��G�r0�
45g��M�0�� [���T	�nx��W��Jgq���7��!b#v��������]�([�8���_�*�;� �q���V��O6��Ҧ���KQ�S��<�Q�\�c�Ӆ`��L�vsk�+��m�����8�T*�Q�T |���_l����Z�(W�9�n����~ƿ�0����5�����x��	�h�]hКdC��"���7�gD:��(Hx�$�C$���9��1� .�/N2llԾ�Z���]��7���С=�����"n
Kg�h5%���p�6���u�h1��].lx0�W	�_�wb�Z	�u�h�Ol�nk�"ϩ9��g��B'�ވ�rs/����F������բ�-J�fuhM�g�Qh�ͬ�tS��N�
A�r�Dc��|J8HDd����3,�!���sWM�CL0�R�7�:6_��R}克�"�� �Z��Lc�2�m��@�X�����Ҳ7�hd���sc�S���1r��2W�Gc.�ߊ�+F����Q#
P�T����J��o�ˬU�Edk-?:r=Y�j�?5Di���V��#0S)�v��߀�J�q]���#I�a3ٺ��Ģ �^�����Ki������ �Ӓ��DPӂD�H�T�-�C;��J��TT����?{�	�^��y	�iRX,yg��b����l��P�R
�L�\��P�v�O~ڳo��Ԕ�K»a�pR[����Wj����0���i�PL;�2�{I��r @�C$nf8�}�������.�6����l��ӻ�B`'�=Sw/��EQ���݈cĵB�R7 |���:Im-����Y�>�:��2=e�(A|;j���{ ��|
�I����FO�Z�1�wM�
�Bd�d�G>�JZ�@(��^G���B�jD�����\���/\ h@��7Ϛ}߄����{�9�5X}'<�~&�k<�m3^�h�f���e.�Y����y�'��'
S$� :�0/7׀n��W���g+^�!S��1�N4~���G��g���S�%�~y�����~���b�L��J��L�kM�8����<�� ���|N���r	(��F�~w:�W�sD��`���~��1QK� Q��S�Kp���N������&���/=�lnlK���S�(_"��r2�c���Da
*^If�6��r���h���<4�
}J�}��7	k�i���y�60= M�.]�1ٯ���|sX�̦�]k6��6۟}��7$2_\f�к�������w�)��09����E�j��46�� �uLn�L�b�v��/���oZ�#)�j�`7�$���>3�s��L㏍<�BP
�!gP-I��'W�������p�д�($���W�����ݜ$(�62���yֳ������%5,U횲%"�'Re��Фq���x:�P�~�T��V�G�������ڨ嘡�K��VR�Z�3��c�S}�Q�W��� �<I�^�����q}z����'n�:'�����ީ<��#��g�mU�{�zp�
�
�5���~e�i���>�e%7���e$W-%,�ʣH��l�B�%��a��h�P}���1g��T0�	N`��V����<��@��gN3I�ykm�,q��,���?���Ⱦ̀M�/%�F��w���%u)�AEdx�$�U6lA�V��b��
�r�D$�e
n���e��<� R�r��%���\8�rDѼ���a��Nօ��1
@�v��C_���aӥ�$��d<G�ʶ9̀7�wR��A��u��(OY�+e��lF�q�l&����{	QP[���>����"
�)��r]���-߱
�j���9�׽��!��������O��©ū�C�#��b�G���1�S&�p���_���81����ĸ�P�-�9�Tw��5��������w���e���r�}��V�O�q)G+��_��	�J� ���~@�KJ��<�5��{簸�X�����װ9�'1�.��ZG4��[��&�4:����
:r��T�?��7�k�go�66����,%[ěX�^	�x���n$E;�V�9##Y�Ϫ�5VN��ׂ�M���r�O�ӆ�x��{�r����&ˈ4耽j���~�����&}���#����(��o�%���-.|OOxG�3��gRV�����.��;:�[�/,�Ϥ���2YOD,�����
P�T~��N�<��h8�0�mi:
J���Λ���Tlϧ?�L��u���U���=�+
lE}�<���ǫa
�D��J�K�2Be��
�F�|��p ��o����vZ���.|i�*�$"��CkPS�q�a�)��pЅ��SgU��wR�����yL���w�2(�=d9�P«�60}�`3��2rts-D��Lӄ�I���~�:n�]�j�� Onϔ=��V�-�2P߂f�vsԱ��J�O����D�Bh�l�6�cp�Qk>�!�%AlO�G�A�5�oh~�����o�C\��lds�Bξ	Gͪ��k�]��Ea�h�g-�?�1Z�9�	6 �yc`��J�3K,�]n�N��)�SfK�)�c+�j慛=.�҂'��ŬR������,k��!�;0a�h��T�H4=��;��E&ѝ(A9��|�q���m+=��~=O���s����N����l0-�^�4(��Z������DF��V�KO���@}�2�&�Ԍ9|�����Lb�D�����v~ӗ��"11k��J�m ����|�n	{���o�h� �B��ʙ����,�>�hn��X7M��bx�_��Vj���D�h���t����W[���/�,�paa0t|`qØI�`]��)�Pz��b ��;������}�h���f������(Y[���z���;�ke���1�8ީ*�,���l�3_4]	�/BG�B�f@ĸL��.��8F3�}�n�z�;��<^��h�	���4��Y��jP�ͱ�G�T��-jtX�閑}����ԭ�n���	�t\�t8���߼�u�n��O��y�����H��J��	ouP֑;�!�uH��kgD���}I}T����q=�5IN��U_ʰ�Iʪ��Jt���K�?w[W�+��c	��98�V9F9�׳�@Yp�,N�|���mN'�{��'�.'�$6spi�*��vr�`��8T���;���?�蒄� Q���>�K����OBs8�R[�Њ�
S�����ݑ�
ʈ
ݗ��M�:tv?�X DV7�J�>�����Aa#��0^Q����5�ޛ��-���:�E8�AY�C��%��Mp���;��!&��}��ꤨ$�t*�DD����OLH�v�LM�d�E ʀ���әT����x'�#�{/Y�rH��0Y�Z1�
;��FL��ф!�P����;D-�H@f�=��&#h�xN�+)������]�<{���7mU���=`�����.i�̦ �����i�o��۳�S���|���������R�&�e�G7��GP'q>�ʹ��xhо�`R�(!>������{j7z�g�-m!��R�h� ��H���q�G�NwY����4���T�f%ϼ�݇��=N@)�S�����)ஊ��UvHO� �{J喜�C!y�\�(�c5u�(EZ��
K�:*a(JS����u>��Am\L�ܜ�-�w��?��Py�Kx�g��k��M�
��fe͇�e��i�A�[��R%�I�*vfW�!�<��^2��x��)Q�^�����d5��k��m�2�&��y( ~����W�Jn�pd��觀8���hV�c*tܗ�@L3���y�Q���aG�j��W[յ�}̋K�_�e�±\1�̿��G��-l�ԣ���+l5�}d�Qd-��W�ñ�^@�0�{���>Ư%��Z�,����?k�sk!΂�Rx8+�����7���e
��8��?e�om?e��e��
ۈ�Y���i�+:��0��L�B[�A��������5ɉ����m?�!(]N�h�4�s��.��y�>�ˁ釐1]��t9i�ap�����<m㑾�D�|��B���w�Hx/m�I��ߵ�M��u����Eİ%|�%kZO_�epi��Dz�e�J�.��`](c`A��p�z�&w��|�K �aڵ�7��ֳh��3XxA��g��V�j����$Ik��JM�u��S���PZ���Ň�9m*s�����ӽO�s��� ���'a�O]u��eЪo��d��|��AYт��A[�\�l������U���i�5X�u<��Jan�gm{���SOp���rAPWuO�?3��NfV�=�@�'B��;YtDm���3ܻhU���V� ęc%�����
����2��.Urz.Эp�7����B����Ip��~�H=�ߝ�	՘��Y�M
b-j��=Af0$N�!�m;�Ǚ�%�|�Cr>L�铙���̸\xN��^�bsw�ZD��J��3ų �V��\Zv�����_J�yXU30-	T��o�}c�*0{��h�bd�(��jxMy��6쐠43�t�����'�O�=
7Q"�R���hi��E�M��F�k(���k�4�5M�5<��M�^�B���rQ2�M=���\W�`��յP ��"��:��[�Xϥݞ�Z��[#��2Qt�'�2�7�P�8���:���X[k�?�r���W$ ��j�p�=K��]=Cm�ʡo�l��㊍�A�0ʑ�Ӷ���sV�u�h�j����x[%����5�Î�:�6�X��[��J��Y`;���mи���NGS�|���C���<'a�֡����3��y؈U2𶌟� �C�L�AT��ɢ��p�/�%!�dt�Do�����U
�\iU����A���x2��>��j�BM��$)wnCJ����������``ao)}�BNՆ�'o�Q��W��b�F~��~� 7k_���_����/� ]�ҳ ���!�ě74��)4������%u �!�4���^72BM���IJ*���_f-}�_)�g�f��I��>�ʏW�0���i]�%K�R�So�� 0SN�,p�Zm1.&���-�aǖt��=�rtG�~�e2�-��"�By�(ϙQ�ܖSJ���Ú�����iLIU�
�4���ϳ��u���V#��(� ���AV����q̨�lq8J�[�ąָO�<*v� �KN����