��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ��%�͉֭�;��B����&Ȅ��n�t��͇�˽��%􈁆-@TOYEX�c^joF����7��/S�+�pI�4jM�e�)����ztѤ�͢dɊk�K��`u@�ďr6����ShU"��p��&��^䞼�#o�]HA	����pEh؆\[Z�R싶C�[ak*z���*R+��t�[��ƻRC|^Ƥ8z���&U�N�ڞXA��<m+�`>U+wp@Dz�Czq�
�./��2U��"۞lF�r�B��&�hiY�<5ΡRo���l��H��4�}�Ӳ��~XH�+��"C�;{��L��n ���j*�����L��$��X��������i��v�3Bk�~���Nx���`�x�_v�b����R��E�\~���wOF�����W�9��º�0��RL��z�Y��[Iv�Rcy��Cx!���@�û8��>��~��]�1��VS( f�����>[��E�
��GoI�J�!�l�`��v�� ��6���b�NM���J�Fɵ�O��v��|�P�h�0+:��BS��}�'Ԡ"S}����`|.?Yl>��x*��C �D�o�{�p��M7nh���E����Т��sg}L��w$���UNܮ��wrN�����G��|B��%�?.m��Ώ|F���8���b�a<����Kuq�'�#骩�A��Qm
)�8Hޠ�����G�;��H�Ty]���o��'���e�Â�y�F�j#J*����e���>��P�(7�N�UT/��U���2S�v�����2$����C�}�Lx��L����v4-�m<T�����wd���_&bT�ȫ5���a���ݵ5	!߷҇s�{g���� O�#��^^b��\w�G����q���KÔHkg��*ɨ$��5�P&�1�
FO�z;�6����I̼�k\g�������E/���8dL��2�ԕ
�իmu��:7ղ�;��Xq�9(%��'������I3��	4�:���p��b8�����&�\_Z���n?��u�|��ȸ!:?���i�Fav.܅ ɨ{�a{Н������>q���C�.@!o��^�P�=�RU��u��^�,a��S��X-0Z��j����O9�|������rA�c�V@�	�X�H�W=3n��i��8b�t3ρ5;Ld�;;ɻ�e�FV�pn�9���bs0���a^p�"y����_��E~NI��W��0�J��KS�Hx�"HP�����n~�ۣXk��3j���Cﳕ����ftB�?���v�Z2�d桯:jv+	}{6�y�
VH�-��K��JCZ@yyݰ���W�g����q>�t�X�jR(.��g�K���)J\`s@�6B�٤�drJ���C'H!;�j�!ϩZIne��<u��oϲ�B����1����¦�WG��/hBe���H�-W�	������
�೅�>T�e�?&�4��<�t�~Y%�":}��ts��š8vLa��OYQ�	J���n���{�C�/��V�� ��3��T&��x�x�Rz@T�~������2`�^����0��(�m(o����Df{���[��]�B��` ��z1��D+��\��5|��`��f%�#a��J7�n�m��9ؔ�\pq�ZP۔�}'~jH�(;+��}��\`�c�Ufj!����2�uc��6©��*�#�����bω��1)B�U�硍�IK�d��&�i�j��ֽ`��ߖ��Z�]-Ӑ��D�����I�paqi=���K��Q��'�p�:^r���8TY(Y�Yq�eT�����Z<���`��E�C����`v�F��2uľ��zvUn{�4\H���2G��(����鱝dX3|��\���:��Bs{pv�M3B5}�dU��;�\\&]��6ie�-z#��(8�P�D�ag�m�G�1�Ъ�H�ox&b�KÉ=H}[��/ˠ�y&H@Ss9��ɧ1�oPI[���54�&�UT��3��fK��/G&�H״�cϝ�"�%�A�t�awM�X�'F��x�^d�2�]dz�2�-�<��A�+�o4��>ƹn���k�+{�H	U�q�;�wC�,�S�vO-���Bt���tuuP�#\a���8�4�_+2<g����0-�
]�?��
�Ϫ�8&����b��e��.�J�]R��U�����KA���̫�=e[����8Gd,�OZ�r0"���hP�\ e黃��p���U�6Өg��nxv�#���!��!��մ���%SH����z}N�_JEDa�.��˂��!��`˛q�3O�����n<��Μ!*-YJ�
�~ÇP�L?�^@9� ~�ץ�� F��
$)��W�%�g?�!�47���O$}Rv`h�ήCHg���}��aXJM|1.��\h���`q��Rr�X(c؀\vݨ��5̆��xJa�����qz�-2&��0��[�k���v���9�C�0�<ъ���ɪo���n�vn+��n|	s�D�>.r�t�g�;#��,��Ҩ��K�Q��I{z6�ˌ�wQ�"jd��_\x��o���iU�⽹q�R�lI��I��^7��L�NL��L<�x�{K�ÿSp�`��kCN�=��r�<�=0�2���<l�]��>���2i>Ĩj�� �{o�t8�B�M�״ܜ.��Z�������./w&��D��=]�,Sf�(�IO���vy�f@@����i�+��G�����D0�ըq�]�Ͷ(ò�T?aOX�#;<­�Ԛ�OFT�Xm�b�Ѳb�L�?�+��^w� K粁������7�,$��P:w�u׏P�>\�{gH]��Α��
[�� -���:V�����r�t.a�����I�'��!TY/�e��%�/jh++�4j��w��>��� r�g�k1o�O�����/E�0@�d�8�-�\PHqߠ8�Tm�h�������j�u\�1�M�+��$�+!44w���q�H=�x�S��|�,�������8���ԼJ�:Ƭ  �̙���m��,��i�k"���=kX�|l+��:�ʚ}�Edh��ר�Xa�I='w�jy�QD��F;���4��0D�$��],8Wlή��:��a[_��w���_�Q�%�MvK$�[�ndwq�;9��p�"$�u����x+T�'�b����O9� R�$�~���W�r,����YN�d�=���lxJ�r|ǯ�5�N+f�Ġ�}g�G��32V�g�Ej�Nd<��x��{�R�C��m8����NӾW�h˓9����E�3�	�f9��@< Q�zb�#���/=�"�������
K�em>ל��1ެ�f2z ���q�G�xp��H����M��e4�������%(ޕ�`i^�?�}����g<� hε��>vA����x:L����^����Z�6�|/:i�\b��j�)�Ы�� �mUr��*S�^l��"����4 ��8�"9�Ds<�'X(,_B�Ӗ��!�n8,cg�!�;������N#��X���?�m-�r�U�#�[d��E���O���=cg�П��h�ݠT��`��ŊU����A
��{�A�ƍ)Z��V�gL4�ܫ?�1�j��������7����v���x,v�M�$��E[K�N-A�>��ݿ���MBe4�%�����B��N�Zq�r�1�Z�
�t��`�c8:���UmT�%�E&*�^Fcڟ{Q����'1�*C�x�踚�1Bl�o�����6�$ÈJ��,��l6I�^np��F��@�䓡�;̣`�� ��Ξ5b�v}R�`5I�
#�*�����I��؎�� )��6�Zj��_�"x�&����g�%�&�	[��w��[�G��%yrb�%ėu�����M^�:&�5�u?�I�6���L�Tr���?G>���o�T�S��#�Z��s,b�n�y�S�y�qiCi�j �qsȔ���MfC�>�.a'�uT���T��vļ�� ��}��7(D��v���߮�����>�x�d���?��A�P�Ns\�-Z��T��"�" ���a���e�znQԈ-�'��5:�#Jx��BD�ӨLk޾���a*'r�G=JJ��_�&��j�Z,+``i�0�n�x����e�fE.E�7-���V=��	�-�7���%����H����o�G���ϒ��Q��ulq�r����O��l��ϕ��5�z��{(�`.M������?�Iv�b�֍�tW}AV�5��e�"��k�A��Y�=�����l����u5��c�ɿ��Wz�f[�"����d(p�RL�r��[��j�6^[���\56�`���7u.��P�r�L�R�`l����&�E����aY�r�!���U<��s�V��G�Rz��:�3���T��T��<j�>?;;�nط�6��V��IǗx>RgC��{�I���2���aD	�m�8�tKN$�9YP��W�͏���S^q��~؟7�t�y+NΧꍻ#����3�P��܉�ڠ�<,~c���[m?�����I�#W�)o<r���~����f@��m���ߝZ�4����Sl���eHdȚ^iǀ���{w1{���K��C�(1�md{`;N��6V�C������ �,}��rwl9bo�K��v4�v6�Ա�*h��1����W�z�s�؍���Ԏ^�a�gHσ�a}��d����WC`dF���t����� ��n�eJ{���[_�xUg�k$�'�O,J7�*�?Sy�)���r���P$��g&��?�����ä�z�0,�3��%�oo'�h}��J���������B81b�����Ӈ(R=wN^f��6|r�(I4|�$#,�i�=YP��IT]w��+阮�nG	�A��U�욕%stn�	X�&h�����Y��4�(����:�K��31�h�1(J,�%K���a�h'�b ���S�U��E�=F	�/:%ν7������Jbߌ���Cq
�YȐ�{��5��N��޺��m�(���Gz��lCٴ�B�{�y�:&��UA
6?�L^a���A��-����X�|�pSˇ�a�H2;�P�߂q�t2_}������# HQ�ܹ6�Wⴄ(#ÊY�RW�6��ڮ�ɢ^�.JqB�/��o��7��^+���Mh(8��w'�FA�s]#�fk�!�a�ŕ��D}&��!e����Դ/���K�>�r���nM���3�F9���4+�b�仪tQ������EW��][�l8�ޤ�d��uH"����K�)H�� ��=Bp�I�%�]-W3�4���fb��#U%k�e�GY	^��NS	Ƚ�A��<�\��l��RCf,�j��'�}n�cR��t��37s���a�q�C0�Yk�@�O*٢y\X�%�ĽJd1Sɩ����k�O`}�G13�f�֢	͖̑�* xJ�4J�N��\�|]�Ȥ!��Y�Qcs���wtvI3�f]��o��K3Vs�x��27�!�i;<����GBkb7�oM��N�7�f�{�v<�'x����|S�n�:��u(���zq�"f��cu�p��(�7�1H
m|���e���l�"5>数�k	A���vR�j�5��#�n�̱���f��?g �)*珒��g�y>����L ��k��5j�E������5uƽ���#A��4P�KE�qb��N�����V4���������3ӷ��G���V�Ĕt,�����Y��}�db��u�2�n7���7?��}�C+~F91���@��R>������G���ϯ6�sg�ۯ�JY9����/�C������K�y��|�9:���ϩ54,�rb���!�ܐl��(�� X�KR�UT!+ꃭN
��1�P{���ܠ�(���_:�XL��V]JR����6�&���;�]٥�{�~���=��	���M|aTᎮ�؊F�N[@A���Xr0�6�v�Z�90u�('��?�g��V݈3���`��ɋ3h�>�挕>k��Z)��Ad��K��z��j��ek���/,�Zq�O��6Z�A��FeP��z�h
�F;���}��`��0)���Z���B��է��e��t�e�;��q�S�7��m�4��k��=�m�me��R�0�����ȩh7$��i�_�")V����� ��+�}]Q-��&��pj����u�fM�l	��2�u�?Va���B8bS�J܃��sD ݹ��ET�P}l��w 1������t1��e��R�iJ��LM٢�<�ydj�h�^��{�̵���+7%5���G[<Jퟶ�������������[R
:t<hh��� ���N-""x�aO����,�<-9g/�Ai</t�pVYEx��x�3���
C�;�Hu	8xM=YL7{%�g�HZ`���ߡ�mM�o���&x�����׽��$�o��$�>���Ø�ҫ����)�OI�u����� �P� ��p�
�&�>����a �����!��3��6��knA�������ЏS��>@���ي��B߉�7p���f��S�o��0�8��Q��{[���-���ʬ�����ְ��t��D�Y�W�5%�07��ϊT����%�a6%��Þ$&�&R�ک���|>F�2����r������	�tx�
���ޱ7��E-�~���5�M�X��]�rc�2�媓��je���2iL�9sq�E��y�d���`���&�j��U��c�� ����:)�dnk�3�G�n������j���,a��b.�M�]�bo��-.�M�=Ф7��@+(�g ?x |�1I{��׉�[�q3��#+̨Yv'�zR�i����*��wA~�ك-�-!PRqE���D�_�%1�YXF>�<����e��|��!�>o̅Ѐ�1��W�AޱR��S��8�����R��"y��iu<��ۃ��5U��Ţ9���R��7��J�O8�ǧ������R�>�\�0�L��$l�b�Sݱ+��F����P�a:o�|����6��	=-�!>�Z�7��;+�ֲ�+P5as2#�۝����fEYX@+hy����u�=E�)ʮl<+�u\dl�UF�Z���t*K!������{��o��p��*��+ŉ�4l<18L?��%�Y�k�'Lx1���� ���k<��s
���9��v�	�����y�J��rZ[�$�p??|֢?��(�P�cv' ��f�yQT���J�5�ԿL��$_*��v
z��U*��A�HX�ٟ� /��>�Az�Ăxʱ�wU��x�d��N Z�`����n�����S��2��*��7;"Ko'钹%��&M�hI�:k�L��;}�f&C�$X�:�>�'�e�2����B��s��Ί� i�b����ћ� ��-c?b����OYQ�/m��`F"� ȷ�}��<�Z�d���)H���B���-<DI֡7�,MY�M�^��*|�b��o�݅)l|g��$J)�����"���L9p���,�6�Ǝے���I�'��\� Bv5Z�z�OʽkT�,s����1�C� u���d����l h'd��:�G�]{1M@�d��O�?� �ۆ=a��հ8�"��o0<��hca�C��sO����W�W4�W������~��~HҸ�_��"�玆�إc�⏫i��K�|�Dz0J���uf�:\�P��;Cܙ�Y����Ճ$ ���>6wH"��.?}3~^��&���i �@5�f�?����g�5��eH4�Y�[�i-����H�h�N!�<M��/2E�=b�49�?��3G}
�<_D����ʺ�5,�0ʎ���h2�T�S�>�<�1B�]�(K�D�8#�I"|�Y�Am���lR��5k�̲Ήg��l�ѓ��P�!�g�A��%�����Q5H��|�_G͆�;\�٘����'��"���t�3ݝ�В�A�-��*$��=�H���\������Ja8�'�1�O8��̏�#i�Y�dr��������0�!�f�'���&�8���p�`8�U�;����k�����n��G[�ٞѦ�h�Y���oz��(jP5��aĉ웳y)<���o�`�M:&`.
>�&�2]�6�4\�f�js�ªئ{���ǹ�!�O���l�U%�0@���:�M���xU�fC-�>.��nj;Vp_�	խ	v�i(�� �9��6�����-ә���-� ץ`���t�C���ю���������N�<��*�]H�E����e����%���7~Zޱ9��k.�gj�P��UGQ���qb���ϋ�z֟��V���Q�_$b�W�@4�Y*k��F��d}2�ڼy7(���\��ߺ��S�3��{�72c��?�^qLf��J&�ɻ`��I��,(�����J���BԻ��)�r���կ�R�(�	����!��[e=�Y���x9��e����D+���7��ݢ)]��e��,d��-�x�~�oa ţ!�M�����Y�0��D��ln%-�
àL䨐Kc��F�Ħ�$������ש���4���x�P��Z�
���1SkA%��8�o��L	�-� H�p��xShq*:�b���6O �8O�Q#���vJ{�3;�+W��|����8����I�HpE!�\��M-�zG�f-hM��4��ל���?���I;������Wt�̼�s�7��&�&���a�ZZ��� puN�i�[?�༏	ո%?H�~Ttwu��`�&�*���������^�#��Q9|���9��F�u�MsD��U���!jZ蕳܃Z{��1�G�ʝO����-4LS�o�PR����D!�i�����_ �eB[�a�)���F`^���r'�S�*%@W�EZ#�QI6�jBLk?+[uU}�tƨ��.v�*�g����w��h�~Q2�`�>(�:v:}����Y�U^�Ox�����!��z��n�ީ5.s����wr9�F�J��A����p<���bVVm��� a �+������Gi���jC�>���ׄ�0.�&�yN�kN�sl�gl������>�uz�7JDF�nM��ˮ��)��$YH���:d1_9�<z�����'a��L�� �I�����;p�ə�W�6�ˤ���\�ȫr/�?}���y�B���I��+��w�
`~�=zJ�I��e's���� 3��,��SS�`�şd��{��2S�9�8x�ۢ{���S�$L���dw���?%h r.����7e,�)�Ԫ��z�Bş�\X{���>�#;]׋��I��N��D�Rdɟ�ћH<[kc}�;�jM�����cR)U�
����#�t�� _��t�EUު��B:/ޮ��Q����"TgȻ,���G��d@�̮��h��x,:����Mz�Sʤ���Ic��<�r�fZ�!,�a!Y��3�L�����z�I쓩a�\d���t�et>.���C�MB��ML����;����ę��EG`yB��]�U͢��^|j��a�?��Q�\֏}��O��p��񭪘Nm��~�H��Aj��&!����ӑ� ��(+^C��,@/ܺ̚E�j���m�^�X���a�ʡDr2�(���7�DU�y��տ1OYp(�.��-�)x��q�Z�р��dE��� ]���u�Є�X8��d  ��6��8�� ��ڌ��в���mY5U�?���y�8�!��^�V���
=��왇?$pq��`Q���;���z@(��<2	/��B;����R@=�s�t�'u!o�E� �A̴�r�U�9&�	�ڿ�,g�pKln����:������y�1���.]}�Ό�m-L��
�-;��'�^44?��ѯ��alC���`�%rhtܱ�N�OM��f�<S�A�����:��Ɍ>4/e#�c�=�����״������?\�щ=?��!��
���D׼[��3�9툜��18�ߞ���ԓFX
�����N>�Z��N������[H��TC����%��e}΍|g�$=	(�8�S�d߷a���ݾ�8L��/��@Q.UG�MMD;B�g*f��_�w�끒��#ph>����:�%t:(�,� �B&Ĭ�(l�x:�4�˅��z3�p�תŷ1��X�E6����| �<�W1�@y���p=��^�H�,N�,s�D5��m�Fl��