module request_ctrl
(
input 				  		 clk,
input 				  		 en,
input                    reset,
output                   ready,
);

endmodule