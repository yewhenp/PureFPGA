��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_���v�;3����ZPGO1<2G���C=f�V+ń���h���Z�|�ƴݐ�V*=7O�t�� �M��3��݃U$�@Άa����)~*��ݓ�R	�RVD�m=��8�AØ�6��|a�I񜲈���.Y�W'�>ՠ����~��U�͇��*~��2q�!D'�rl����YF��'S���W�G�����c�s��SC��MQ��F�xV��n.��~�V��$fi_�i�P�D�%_�K6�^Z~�+,ˀ���b! EB#���Sc䐎F����VIͅ�`�N�Zl�i���I��gq�|H��c6�ٓ�[/
vl���N�A6۾H�sűdE�b���_,]��6�ö3����c�Yej��y޽Z�X!�t��53}0�r�V��2���(X�y���*��2�
@Âш+@��RnT@�#�^������W"�˥�Hз�Lv��F[]Vxx%]�1�LP���ę����yȡ�k7�nԸ�x����nM��ٟ��K�2�(�'`U#�p{�`p���܊�'�*�0[�W��o�	�4����B�E�$���5��f*x�6�m`4q�"�!.v ��\7U4����3��O:rA�8�����s)��2S"U6^+�o.�,�S�U<�~�nm)1���Ɛ4��-���Z�zԊ�p���'�Ek=ˠ��-K6b��c�k�kvp�ڛ�G%�}�F�j�P�t�=-Oꮸ�1ٴqeLƀ���wÏ$#�F�KS���S/������9:ǟ ��`E��=���Q�k����bu�8ky��e��xd�_!���K^�QYʾ�$Q�u��r�fy}�9C
Յ~��S%�]4�^�%�WA�"�����I��[�\�SVM!I�w��m2)\Ӡ`����F#��[�l��,��KY-1�|w� �E(@el���"D�`J�>�`wǫ�Ɂ�L� ��,d�	�P:�O�0�
S���j
>�T�RwY\�T6Ǆ�	����S�ׄ����c�G�:�Ip-)?NA�Ŝ��Oe�D�]�d��`_�WR(�^���˾�@�
xxW�6��r��S	MM�t�N�j�'dӇ
%��p���ښ�����t���gۜ��1�9Я]��,7�k�H1��n���ZmJ,fr�~�����(�)|�:����F����+m�Յ�N3�,������%7=�I��g��LD��)qM����A^��M�>,���;�;�Qrc)K 'u]���!�é�Z�[Lf��)�#�B��SC�aћ�Wz�'�AM�⭁7Q�@��N���rH��UÚJ���|��p��C+Υ꾭��+,T��X�P�^��+K�3�qrH��R)$���=eIX�IK�N��LY������X��'��So�d1f�6"��k��kR؋�.!r�Y�BƊ� n
k�g(����	]��C�LL��߽�Z�ݿ>t�Ǔ @tt@�������sc�0-,�R��H����d/O9"S�	}&6b�Y�)͈�����Q�n�)^�_�ox�f��̉�˚�3f��e=�RN�y�YY�KT�"^���}�DW�T[��ɂD��JW(10��W��(�!��I�w1_���������F��eIs��"�WaQ*�]��!��_���i��6a
�i����⣈��,D���(䝭����Ϟ�z�-�����ה�5�IKZ�_I��@YUz���֘�uCc��C�t ㍙3��/��4��p��Y�ǩ�e���>����?�q?���{M�;��m2������h�-XٽA6��&Z]�
�So�$�1"Q�b���-��cjV����|�֟:��c�F��Oȷ��|d���	��Nb�kp��E��p����8�V�#b� ����|&D����+�F|{<q��Fn	o�ҟT5���z�i��b~F�f"2��孳7b�L�Đ���w�����b�|�����Ɩ��?�qg.��������î��_�C �=N�.��8����אlb�Q��Ń<�@/��]����_��N�@�0TÍ�VӐUo��H�5X����G��L��Q���N0�xV|�?��_g-�FN���I�e1���Z��vI�mi�3_���	+�ޓ���Q��'���G�|���@̶�%Q��$W^R΁�k#�V�Q<���G����{P�7�I	��4#����;�u2Zo��Hts�O���U�f�-�:#�v�����)o���.�+��Je��K���J���꫆�C�L��~�0qB+>t��'�F��3�b&/#�2�G]�4R�?��Y�P����L\d��&���s�����q��̏|*˂z�n���gF�;W=���N��AyW�c#��Q��K!�3��wT�KP�w�Z�Q�N`�@��{��@���հ���,��0�W���Th*�t�:�8,��4l�Q������b����*_ciL�j7 �I�8M����}�"�<u>"#�����^k�]�=HJ�f�Ϧe漉W�KwJ�}�a��@tm��tTg?�E�����L�l9E\}���U�Mk`�RND]��D��q��U$�2ܟ�m���p詃��������_�w�R��I�U����1�^��n��Q�R3%�E�5U�5v����솫����I}�%�W��r}�g+��?�?���k2%��/硊�:T�D�:Il�Bq�,�Iy�7�RI�f������'�E�Oa��/�W�b]�mU�`īW��L{=�h�?���l�'�m)�}t�A��V�r���C�BX\��ٸ�%�K��+(18���[/(���C���8��W��$i���Q��Z�z�V��-��9ݚl��u������8&����Dr�$���Jf��-~�@<�f0g����ؽ�7��X�e0� �9��G�L�qJƕֶ���^R9�|d7˙ ')����L+���_3�����M����������1[´f������*&��XoZ�ل���-�ӄ�Ւ�6ՔD�gq;� ���*��w���ӿE��y�紐`���W�[J�w�al��e�~qq�%!�����C��`�S<����_/:��Cy|�Z�c"��$�����K,dt���$��T����d2�ǘ�i�u�}��e�����7s��mK�H�)i���(�&OS�	{j��L#Z���G��{qK( ��^w��0K��{T���m�(	|:5�3�q�H�a�>0�fsnHU1f��%�@��z��<>��������̵�/��6c7&�U/��e�kٻ<z��!�_1aj&�(k�w�O�U�A6Ö0��@��[���7
Y�kQH�� �>穏�m��]�R����A?��o�1#2<.��@嚩�=��l8� Ǘ�}�h��$4�&�6v�E�fm����	+���n\�f��"�6�j'm��˸��R��e�hLG�˿sPD�!!c��;��`�{$K��q"�-^V�'Q?q�J5��
_���z.����kb
7y��0	�bѲ������ ��P�7Y7� uI@�!��M�(�Ch���-��,��3p�}D��MY���9ɨ+��$�[�@� G,��������'�6�!݀6�H-^�25�+���}�����2�L��w+I��O�I'���LO�WLw����uN��l4�����>���E�����	�[����C�2���N�[�&�~c��_�S�	��Gb�M#RY�s$gۆO��_���TE��>2�&�lL�8e1�`"j��=H��Uav�xMuI^*�(:��YX��v��B�Wd��J6P�(��rc�+�>	
���U9��({�.�^l6�����y.�a����,�	m���OB�\��� 0Ǖ�[����IR�>�|����ܔs|�{.QjA����қAH��o?�2�6���V��/��z�?r�N�f���U���<RTʎ'峂٠{Bv�������dY�xX��G��n�DR�ގ�@��m��jrN��'�t��*˂�o>�&`�����^@�mW+}�������8�$9��E�= 7���T�e\�?�RgW��n��|��sm8j�e�q�:1U&��)��+:!�^� W'����ʩ�X��B�U�#a�ϟS�`�+��������D�[ӽ�ɖlab˓#K���/#�����"p,��2��Ɵ~M�|�|U�������4ِ�h\0�����O/�������<��ɾ��y���w�T��7].7t�Y��0F
Q b=�F{֙�tc�fk����4iܩ��s�==�9)��f!|D�6S�<�US���������ͻ�s�MGL�t�碨fr�q'e�(F;F�ć�1=<�4ݶ���wk7��%@P|�p�Q� $�~�=�z�|%ld�CmG�l�5�|C%ss��a�|�Cq��ݰG��f����P�@ϗHfk�Y�>_�����ib�	�vN�FlgY#�On ��|0{%�m�<3��NA�(��a�oM��˵�|�u�K�Tj�>c=W���}M���d��캅䮯��k��m�%���`��t���W��6�G7>|�~��Z�N�q�I�
aPt�B�X��K��e؏�{7���!������o�99�w����;�߁��p"�i2��Ȯ�QA��_	��t�J�Y�QmvB$�:XH��X��B��3P\�%H*�����(`D��^	]l)���lV#!�I&B�WdO<���׫��sh��|�ɼ��[�w�O2΍A;n�S(�Nr�K�}�CtzC�Z^���w��"���bE�ǝֈYv"T�<���z��If���,&�l��BvE�@)Xޡn�BGGI��� Zi2݊濝�T6ۄI�Cδ\�d�$�w���d.5Cy�+�F�of>"*�Js�m���#UaӐI�=�,�[��4F��bX�GJa`�_��;�o��|F��y,�"���QY�=�1D�l�MO2��LKeB�(L�4��	R[�Q���s1��C��J^^���Vm��b��CK���D®4��(�,�[ l��J��h*lV5���\�&leOQhQ�ޑ�J����� �&)#t\b\�a�׮���*f��Q��1jG��^v����x���0c�{%�������R�Ix\����ǜ/��5瞇��i��8.~7��ͪ�ת�����*ۊ;~BĆ���{]��s�2�5��^a����*�ґ'*��b���prFD6A�;q� �2W�6�w{��<�B�>����y�͝� ��V���'���,�8�B~d6��J�����2�H^v7Z=��ʋ(r��Pc=���Ӧ�ܩR�)	PS��kU8!^ᒕ}��0��2� ���bOUI�k^J��)�!�}m!�6^�t��H"�=�5��vl�����y��
�X�jg�����t�=�+z�J)<���-3�Op�HV�����4�B���͵��������Ɋ�
!�k��D���� rF�*�*�
u�C�[���EY�;�[�[�]^���J��6�S�W>DV� !��%FMjΟo�є��K�� qx<�����I��yK����{�g@T*�����Jh=��X'�X�.�0>f�,��ǀc��-_��d�X@��^���c�8'�mw�����y���:�"����"fEQ����E�H�Ҧ��x�N�{��*���H$� X�lI�������&ػ/�ڭ���W7��-6��]�pϲ'��f]�1M�b����1�m���"�@I"U!j�}A�4E�y��nl:?�[� ��n*џu"k	+u�SH�.�zr,�+�C?X���7F�V̵�	+��D��p�)�E3=�FJ�PՃ�S�>k��v�V�3�km|�����2�~����[��+�y6��&#�|o�YRL۱�Z��ǭ	+[cVɆ���[��R�(��@��o��PIn��ɰ���מ.Qm�݅��I��R\����
т�I)Q�]��i��^��$!2���h�HK(ϾT�بD!���Ё��*�