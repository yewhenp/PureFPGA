��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_'�s-�`��f�>}�V���wJ��3�o�ۇ��.�JP6�7��I]|���PN��uI�J$ng`��3�y���0���zL�"�i����������.�GC��V�?�r3yR��3���_����O\�WJiq�W~�u/I,�@H�>;U�����0�Y`��s;�a}T�Z>
*
�9�>�g�J�mD���H�����|rAN{t���1��g�m�{J��1���W�a� :�彶`	�lY@0�a��� �u�|I3��uȅ�:2�o�K��8m<x������l�Gu)wB��M�\N�:�� e�S �H���`۟�Z�Z�WI���ަ�Wo�
e�	�wg�^Y��|�B��?8F����,���M��W� ����˾����V��="�~{a%{.%��y��S*i�-F�w�("y+��-�cl����4��Խ@O����\��7�����m�DGP&0�Ǔ/̹�J�ߪU:�Ԡܶ�����|7�dA݅L��)Y&�exj/~�
�?���1�.���lLV��byłhOG����'Q�q��#
y9E��c5~~$�H�L�a��NU@�2������1�r9-����JBwb�/c�������'��c�yH#�J��Y�������̢��_�o�ُ����;�Z���<���r�_[>�g�T��?2�
��#�������I����!�k�^0�.�,���88$�q��/�oM	Y_��5�t.-�jL[�Yi���C>5����>�<��̋L����E���:�3�������7Ts�mȡ�����+�!�����>��*��� r���5(å�r��ΐd
��R��jO�X�'�q<����̔��cBq�)�)DꌜJ`f�!��~��mg/�{��D����������@dS�)�@�W�eڎRN��Բ����`C�����[��r�8�я�y��I�@�*�r���ܠ����x ��SC�M�6�-Z<R a��/�Q�vj0W��2\���S�&Z'��I/��L��0K���O]+|R�dTӏ��� �������:K�"fb%ta�����L���Ǧ�h1"���9`�=t��2�������'N2.�g�Tp����Ii?I�ļ�<G�5�r_.mI��ʢ���r�+�YpBv�����bmcz��V����*x�_�T�CB��E�9� 9�.d���2�5�$ð�eY%�-���|n���o'�h >��S����:N���N3&ʢ�h�O}��� �@$�`	�=���Qa���5cb��G#��*�	�20�E�2��e\�NA�R�X߿T�`���#i���?H��ƀ^_�gQ&��7������&)#����`�J�H�7uk�eۺ/����"|�|�Nt������$�kS,Nx_��?�ppAQ�+�+�b9��w�f�|�-H�t���Ȯ͠Œ�Վ"@����U�uB6�=uu���&֏]����,x���d���%�&vTDf��o$pY1��y}�K	�h-�������������R�F;�?夸���93�S}�E(�y�f"0s#:I��#��˘݃(+�����}ρ>�/�/�7���)=بp���M��F��U��S��P�)�(���H����_�;.@vE�(H�W�0���	�^3��B����,�}���{.�\|5�4MsL@��{�,C"2A�Ĝ�1�G����Iz��T)��:���f8Pd< OM�i�Dp�Hm��fj���O����&���+�+�K���Ml^[�Eyk#��	��]82#�����<,4c`#MP�6��߼�ݵ�q��C�:�J�r�4�	���$`9|GQ��Ryl0�kp�C��=z+��m�aL�&�b��%k¨ .��+t]�A��3Y�ݮ�E�P����t�aU�՛�3)�f��4���$�g��]�5���-k-��tߺ�QwT5��Q���Ax�{���!��,���%����2��Ҙ\��r������<%+� ��x̝�,�V�K��J��=���Zwq��r��x1��]�>؅���#�&,����t���I3�-qy=N���7Ab<O��Wu4X��1��%\|d�w�o2�^~MU�Ls��`�f��Xqk�lYr�'[�W�&?}��!����ꟹ�sk�dǄ���5'x0���<�q4u���A��:��k^�!閭r�72{{���9�T�h?�B��-6V�J�>fB,!d�A`�C� û'�I>��;Mʐ�Lv��Ӄ��*��ޔ�! \�)Iv"�¯B�	�/9������A����7P/����4��=��Vp	;��Ϛ���d)�+rO��%�#��蝤���&R7�	���+��.��5���\wG���m2g��+������Iв�D�×�3� \�\����$���/��:I`� u��VQ����	�@ge⫙��H��oP�|��f��|a�s,�l}$`V|Nv��s�L�h��b�$H?��ew��B�J2|� �p��1�e�>*��O� j�N�z�aoȢ-���*3������DPi��y|���g�~�lv�����_�s%����~M�"���.�h�ݾ~2�S{��}�N:T��"^ْև��?FV0���L�MKx�Qh	��)���:WQ�hWP�%�����̄ڂ�w��;��ϓC��k�X.�v��@�qL���I�?i�T8t�TuEzGүa����^=]y)�4{�كЩs��'pN��%���Cc�ٵ?�:�*x� 4�m���3�������ճR�-�L��52��t���,�˲����sT+���]��B	��ӫ��v�����rp;�g�fdH`��D���D���Xz��y���CG�|ޙ�&���R7�a�Ib��`����R�)\�_��AsxKL��@�U�
@�j\��%��D��9���>Ab��J�,!�h�S�~�Wj^E���b�3JS_�X�"�� \#%1��E�bń������.��G�҆`��L��اs�xW���`�`�4�F��y���45���;���';Dn50H�~���`��e�&R@a�KH)�N��x���"�ͩ�6�ҋb�1��>NY{�-�1[�Y/�ՠ�x*�T�/�)�_rO<U�=�Q�@J��y�}/C��t*�!�u�_ݹ8�C�Z��C
�fbk��𓁁s|	�7ru�D�N4���?�=�i��~�>�-ؒ*��m�fN��٦f����8��}PW�yb�.������V�b�h��Zy��g�l����FXC�^�i���Q�70`�71��H�׏�m���,�%j]�y��[2x��4ʙ֥@��mSm����HUz���*LƆN�P�)�2�p�+�"��z�_� ;��w���ƕ��<U*e�tO��\ð���D0^%�WJ+�5�B�+sկ߳������y~�:��4��&`"�",݈�
�X�?��[M�9פ_`?��Dr���I�A�� �}�r��m1T����(�v{pF�^5���O�
��.)��Q��1t"|��� &���'�A�W��a8�r�A��Rc�p|a�y�G:� �,s�p�`�/���\�Ql-������Y��!"0p{ī;wh-��#3{p9gY���vo���ҿ�@�������=xA��"�*�$ԇ.Xm_�������P|����7���C/�1�@�g�m��*W�֟��2O�|2�N���|t��2<F�
 l�z�|�*6�x�&�o�<X"v	B��_?�ݎH�tL��w�/�~�<�����ī#�m�C�r�F$���#:x�y�g^���E�P�_/x�.�*���m�������J��C|0��v]&X߈�wZ}Ȣk�bo�2Ց:��Eх�_�$TX�h03T�3���@�C�ܚ�p��%7�?�)��_�}/����	27��7L��$tIܤ�.�oÇv	� ��?�3�H��>¶�Z(���|��P�ogt�`�.)��GK���P�ͳ�Zr��?�4̑��7ƭ�����.3�� ���K��	T�Z���6�v@����$,}6���Dt���}E�<A�����;�LS�݀&Qx�n0Oa<G�1�mN���n��H�z�4��yP�o���%�'ړ����U��c�̼d��|�MH+��#jSҝ���s
E���kX�Kpxw�#M�gU&T\�#��ѧHlά�J�4��̬���\��)#�&�8PY�ꗂ�����[s�Bt�7���i��kR�0�8� M��	T�?t}�S�]�O�#�䰊�:A\���1��e�L������y����mʒ������Y�$�(W�2��e�0��{]�Ԥ�.���S���œ�'^�j=
V�_.\��?6��(re}��=����v)҆3*`�AA��;���Ж�,�SpJ�jZ^�a��gе���\>-��!��z�Za(�_�:�4��Ljw��v+Bgي]P�
�K���U���x�䁸�Ŵ֤���>;R,�dC��W�k��r���z�}�U*J�&I�����WSv�zRy�):���,͗�Ñp�q�����5R49s�F��qM����S����"�
K��ֽ��ʶP�� �N�Ayӿ�|^�E��v�����^���c��X�{,�8	�G��"�E���5P?���uA�,"T��NB�����V��4�#�a�O_���=[���U�d�M/�p�����D�y�9�7S�0�pO�?��)(Qx�g��	���0@�X��1���}S9�R�������浞�}��u��m��PK:��&Hq1ӔWԗ'�Iƞ���h�V9�ʰ�7�v�E����Z���G%��4n�Tf���E�Ǩ�)-����E��_�ǝgFba\PY�%�iɻ����=[�r]V�[<5��^l����hm�K�@�����L��]���czn>�׭n����3�&&���LV�G��a�f��	�	(��ju��e�B*�g2�~�3�\���4k�t���5������uv*��i9vۢ��QOd��)�(��&�展�&'��ZwYF��!�i�P�����*��r#�ޯ9BOQ�.�-�#I��WւB.���ܷY�nw�N���nHȗ�*2Ӧ�z%�5"`�Q	�d`�
V������)��v}$���m��/�Z���<���d�Ҳ̟�H�+6Ê�	z��P&��aINuk��\���n��e(_֒��o��N]�$�(,��yA$ϕ3�!��I@�mB"�a�3���*R2�f���`��G�fO]_���$�`'7��nK�[��*x��IH[G�	��UP*���F��/#T��ϪV�'��*au���F�c��7[��M��QN�qOE{OB-Ø���[�c���ŉ)�1ݚ.��	��۟����<��S�*{=e�6���+(�GN��O�V/�TU�I��N�8��3)�1�Fղ C�%�D���{�;&4߾��rT��y�[�V��k
 �m]:�����D3�L?^~�u�;[Y�FWL䞙S��(�
������=H7;�\��8����e�ŋP��?�T���#�[hSt�B�h�G�`��:�?ƅ�H��kz��<_-ȭ��[�b�g���CKbacBt8?I���cos�� _����ֵ}�:~.�Ua "ߘ3(�l)H��]O�(;��Wf�l�B�b�,Z4f
7\��R�u��!3Ôk��G�uB'�WU�OE%�Y��p�d"9��;ڤ���j�n�yl��Qɬ��RBR�t5v~���=I�]�z�zh'>f���S���#ڛ��ʾ)�j��Q��~1h����c�������6D������"���{/jF{�2����0p�Z"��W&���R�}�a�Բ�d�}��惛L�����N��|��ȄW�je�OG�7�
g���TW|bzr��m�eNӻ	�.w5=��\���`J��{�§��n�ehI�z#*�����v+y�喔 \��5=4^4ʭOi�;C=B�c	�"R�C�BmԨ0�+H&&'&ab9��y{ik 9d5�Nh���A�{��
��B�
k����6�,q+��:�I��q6������֡.��<�P�Ʒu,���g��s�gc��uY��j��JG)n|���5-~+x��L�!Avmi����ܠ?*}1X]`�ox{l`df��[?�x��_Y.,F���OÒ�u*�lZL��2RT�>+�&���Z���"I5������!4�pm�n�'��L�i��u}�f	�%��}g^lp��6���*��4BN�oX�����Y�k�W�G_�:ݚ�rh�Z�+�Gx��/k � �S����@�!%.�G��˩�[5��'��[*0������� l�v���Y;�t�3�g��"4"�8a�j���P��n�ZOa[8h���i%�܀�������?�Qn�M+󈐮�b�p���N_�N�a���xrK��?�$�(��gJ�,�kjH&�+e��!�ы"
"��T���f��!�ϭ��>���aU�����}}��7�'��0Ęݒe���s��8�(�O�|��;Ƥ~#BD�����K�=2�#�~� ��c@�s���]/8�[��8�dS�)r_V�>���N��������u�"���z�;M6_X���R�F���9u-�ho�8w�@1ب2�6��X&�@�Q���|֐��H5D�ʴGB	}m�F��]Yڞ�M�V.y����F��mG!��3i�]mi�w%�g�A�����TٕM��ց'Դ�C��(���"����������H����#WV!1Ї�[=/d���X����<	���5�,BH�l���vmtp�UFK^�߬r��$I_'�@�No�g|ٯg�J8�x��kk'�1{�Z��	��x�#��s�(l�dHEI�.-���v��tG/�16���j��EApN.9�&��5D����ڛ%�JE����l	tr��v&D���`��rZ���	zj�J'�;��e����I,M���x�K�mF���W�Pq)ũ&�Bkr�Bq舠*�:����3tTvN��N��n��g�R��ҵs��ӧ����-2��Z�q���Z`��d���9��ۇ�B,����JH����j�����[Ww�����Pw���r' ���#�D�'X�s�Ǽ0����9�V�?�/�L9a�6�v`�k�P{�=��x �v0(@$z��,�c ���s琰%�,�}sM���YKe�ʞD@���Fv�9�To��68xQ�͜�$!����;H��l�=s����R�,�JH@�Ӟ�A�R,!W�����y�Dh��g$��j�'���:����ydl}B����>!~��z�5lݴB�L?�<&����Vp��q���u:4��L�E�/j���٠�	�O�0�K���g����$�4~�{ $��慲�R���n�$ٺ�T�j�P��m|��p��;d<�Z�X't��k0lطm���̿i��c>�Ϋz7XI���p`�͑KCda4/9P6����1q�Ld�VhI��2��^6�>��:Ҍ���?x�"4H��o�"2b��D��BSg�^׍.n�ݝ�'�:�;�v��Y�kY6�2������T;��/�N�e?�|�G�P��x�Guw��X*	��#��+�Lr�$4�8��R�8 §�=D]z�N����	���e�q�p��]��6
5`���^��ɎǦ��z�����Ɗ~�`��O�]w;�����oK����'�c2`%��&��Ƶ���
&h5%ЉdR,�_JZ8?�;T�5����Г�رh`L �����M8��� �N.�KD?0Ԟ���NB6C�o\��¿�,>�!u6Kx��@f��C�Y�M0 ���u���~Tl�ar�	��SN�����wz"�ӻf�lK�
� �*e*�&���l�}�>�*�g���~��_$u�U1���˟��<�� ]1�״��^Jz=PUJ�a_E���38 ?;�3=���% 91�μ���%�#��1�3��H�����4r�rϸ��iy]4u�?�j׀"��,>=�o�4oj3�!+8����b��"4%���u���c���d��G#MbJ��*B�غ����2�*bd�9맼��8/f����]��1��'��+�f����>^��G�����Z4�@�����=�
Mq����ܰ�e��C/�%S�jږ�S1�A_j|E��N3W�ͯƾ�r`��DS�"d�vl��`n=6�ܠh��\���4�}�����Xy��4o0᫣�;=��+�SKꚇ2>��2�6���HD�A���%�&ƟͶ��E�`
�L0���Y��6�z�� _r��.��8U�q�~���yMl
(�	H�Z:�B�( >V�4���m��cJ�:{I'j�.��;�h6Ȫ�L�t�������?K��w�C��a�V���d�Umy�\ �aL�6�����M顢K���O8m�M�Nh^Jvlss(ni���b�n�`h�!uI��o���\��f�ꌛ�)��
���W?�Y3k�֬Y���f�K�����~8(��D��l-L�iK���T�CJAz7��z!-��kg{7����'��W��;䟢͕�+:�=�͎�f�7�y��K>�;P�+��KRT6m��ܽed��S2��� 9�tw$TW=;RO^���*r�z�L����$�Hl[�o�b��dǾa-�8eI}Ԭ{�<X�-�����֚�~���J��Q-�%{�?��;����Rј��MjZ�����*nP��4������زd��nh군=�)-���r���Wr�&�"K���Y�+�.b�jFԏ��B���;;R�a�}Je�^{n���%�j���p\�7|h9xm6<�#�Ө=n:����rI��
C��e�鉎|���e%�g��eb�7E3���xp��Q�J���I�W
�L��=�0p�ƍ!�"&1��x�\������s>�,�Y �@s�a��2��B��l�H�����VW_f������,�&ю��C롯�pv�yF[�½pg}~ӌWRMs�L��->Rx!�CZ�Ӹ7_�/�k�s"�p&�L������X9��XLf � �3��@���ew����GTj�#{�������x���L�5A�n��>��Ŀ�����md��#�h�q�Ǆ�Wo���i�Q���G��s	����gG�%�w�:ٙ��ygB�t�D�?�&GTl��zǬ����QН��{=��d����<>���c��$Pv��[���ز��t�wx~}&���/<�C���%tb��}G;;
�rk�Y����~���
��N�74X�J�$S̏RU��HŖ$��&Q�n��'F:��dd�e�������Lf�"��������H����K�fpj�6.{7ԭ��e�ܞQ��^֡r^R��K��	"��m�q=�s{��{Xa��ؓ�8����<yIR���48֝�aɀ�?P¸ 77���;�$ߘ#�4�5�_UȺ��5�����|�����TB�F��[[D��x�Hw���RY��ܲ��n�m1_��\)�������	\1�_�����<4��e/�gA�~�>��ߒ>5.��2 �u�yd�� �qP@�ҽA�i0[�Sf�T+�id�]�G������%X?6�E&Mݿl�?�|��L3YfK��#qk�7bS����=�w��T#���`9P� �ʉbR��%Mw������P�"R��\y�神FN� S�1�b\����"����,I]Y,w��]M�m�g�!���Gʢ�� ��>-*ѻ�%p�����OVwn���`�΃1�ROF�����'��B��c(���UgN��9>����%b� ��g�����y��'��x�H�o�}��<Jj��[��hG#��I�閻�)�8�߲h�G�%8~�%F�6Y���K�=�Oh��2�b�죰� .G��.J�( �k@^(�y����w5fH���1��p���F�����G�Š-c�	>6$ӠL<<ԝF>.�
��=�L�*!�-�F��<�Hl{�|N�=���
}�oK���p0�'=�I࿬JI|�����g�j[�Mzb��WǍ����b�x�-��s�ߪ�&8F9���bt�+3ʷ=�$�d��ȻC��Of?�ٸP���� K�H�X�����ֹ/�BȈP�}"�d0� �~f�� #Ӈ2�7�zz?��ׂ`L�4.������p��6_f��:����1V@���� �$�Q��8�D���Խ�'g�n̝����)�D�gnq�2�?���3�ZIRl$7}F�j����.�<|�R�wOF��TP���C���Wp�s�a�"���!�[�6����&�P �z"'�=����8t��J�c�4����a�D,t$ۥ��	Ș��A��y�ޮ�a8bG6f,�K��і����!����	gh��w���VES���z�
�^�,���c�+L鍢"�o|����h�6}��6�b�k���&�7?��b`%�!����M�#\��?�Ojlo�W���˥���A��M�?��i_{GY6���qyC^�yq�h8h��v�`+:&��=���� ܒI��yڏǩ܇0�����X�����ے.���Y3��E�^���F�W;��$�X�<&!D_Ȼ��4K��o|�'Ǵ��l�bᏯP'�Z��e{	͎G ݾ�o��EeH/ֲ"?e��T7��x'l�~�����0��G��ثB{K�V����
�5�̂}��g�*�/�$I&.G��L�D�
1�BE.�n��CS�k��!�����UbX�����O.g���	��S���%x� r����I0C[�W��=S�֌���A����R�����M�5�ڻ���Y���GHj���\�,�F�39O�7kߙ����4.
��h�מ<9&/ow��3S���K��f�4?(���7@RZ�N�!6�=\�v@?q�s;7T�aS��4�o*��Ôl*L"�pb,I��2*�E\��"q��݉<���]�� �����-߶�Y.α��ԗ}5=��(b�[���TDK���-)x�!w3�\�
>�d���^�J��:�֟U�f��;��@_O!(�����U����x�n�/cm�a�X��ğ�}K@��rc��
�4�T笵��c�k�ہ3���ўХb���4��J)"֋�^��]e���+����Y��2�0��d-Ⳑ1�������6�#w���5Ղ-�j��r�;b�A݋�b\>.�&�bA�|~O3�H����]��]0�ƀ�3�l����P��l"ia�C�T/Br&�W�s�"�/DQ��a���w�W���n_ɩ,$|�I��t��q}��W�ӡ}k���q@U�N�fco�϶��AC��QP�T?b	�be�nq�V)2���,$O�a�y�!ɕ؊"f�7�5~���Eꗐ�3���4E8�~\ŕ�#v�4�@ g#�X��;�}4jYm�Obt�����+��\�$���G�8�<���#�}�(���I��E�e)F�9\������u`��%�6y��U;L����%2%n�T?$�L�
G(�		dǠڃ�;`���/�$��`�a�q���	�g[��_d��Le��k�"��f\��j�����9�jw�7�&��ğ�db1�`S�v�$x5RlH܅���F��.x0������j<8"����d6�4���.�P:ÙB�g��%Jd�E�5���˯���A�9�'9�A���5A,��~uyaIH�tg���*�%raEZ���­51�YfO1=�%����E�1��gfx�l��1y�uQS���: |�m�V ���e��2��$\6�C�e9�0.Q`�[D�۴.�f�Ye���8��H;����gn�]��dH	���j���P!B�m��xp\S3��y_�$�T�[��Ñ1E/�_<D��~;7�ԇ�pF4�����I������ə�P�p�z�:)�C^&ĄNk�9�u�eI�K,<�FH�֢#�4~��,t'��ܽ�aA��,��nX��#�����}���G3kۣ̽��)[���%�M��r�"N\��N�$�sa<�����`�ʹ(%����ӿ���Z'2-+��Jv�؁�,D�v>��I��i�z����6��Q^(e@p�bY2�1��*,��^A�خ<�!�|0��\�iB�@A�ahoT)���I2d���ᔢ_7R⓬{GvV�OO��Z?��?��A��P;6����<�ß�O�����p�p�o���\�R:���������bB@���%�s���;�/ !4�ŹWm�S���H�x$F�J\�X��PD�}5��"������"žQ�Th���XCE����%�H*?�(��T	w�)����Z>�N{Y`+�%�R7֕��%��Ļ�-�'��E#��X	��k��z���+	�����QzO��b��j�eF}�mj^'�ʥ�Bj�'ߧ�c6��*FXZ�еH],����t�Ͼ˜rY�j1T�L�W�<pI����0 ����X��a8�v|ݕ�����)>�i��F���J��_�=^ӓ�1ߌ��qG	�S��B|�CMρB�����*��V�M�Jl�hC`������Y:�$K��6#��/��b�o �d0�YXY�I��nr���<��H �xB���v/���F1k��V3b����x�hN=fT�6�t�ϵp�Kڕ���"�@x�~}6���/3]��ݫf��y~�����\�B&�]�Tn��� 5v��.r���쉋��X݄�K5;n�~K�%��� ���W����+ʓ[�w��/dg�ę@�)��c��$�����q|�p�>��\�׺��A�r[zU1r���@%�*P^2��Xb�x�v��X$+_�O�wY`.��`��b\<<2b��[30�������^���yZ
W�S*u�3��� ��$uUsaT��x�^-�u�Eq"-��R��/'{�PA��t�$�cm]�/�VM[��}����8%�������n@��[_���sI'�����lݬ�������{�c短�LK�e�������s<�o>Q�[�d@R�1 Gd�X���I�Dv}g��ևlz�5ĺy�W"R�$I������ �� ��n��s0��4V`����z�����{]��	�5 �!����2��kA�с���\��A?<�5wp(����u<lϼ���_۴�Tѿ���9�G�*�=�9�%1��d�:;�g�J1Y�R�g�诌Y|�/q/R�x���Ӫ�!����c��\�mꊣ����%藾[�~����.>���s�!��"W��p��S�/��9\�6�q��t0�=����=J�4�FCrky[b�e�����2�������oRYz�l�<
9A�������w?�ߥU���6�7�b�VL�9Y1�oO�X�?OR���J�mN�+U�I]��L��i	�i�ZnLv`"UY_B{0��I0���G/������o�v^��z^0�6�Ij��|L����K(}�!s��r�a�~�|?`�L��:a'�64�n�	����-����H#�XJ�,K�n���2�%I}2)�>.�T�ž��4g'�#��%��{��S�=�9_e��(�Pa��.���plyq"C}��v���5��F#C�5+UΣ";r�+E"�/��a��.��g5��:�tW��Z���a;�2[We�S?+�`WL�$�#<�X7�l��ͭe���}�~�pI���̚8ٽ�-%"'�d�b���ÒJ��1�W?����g6��¶&-�zi,r�a�P:��?��7h��8�^9[�rn���@�j،�b�y=����]�R�W�`9�E2܏)�aV �?�w�xY����,V~�XWe�!fC��_i0[�+��B�O@;Į��2{&�{���b�=�uc��*q_|��d���������v��� ��$�!�ٳsRסb��<��>��w�a���J-U������1�s;"#�XT�����&�Y�X����I�����`����!�0>m)C�%C�<6�'ɆBk��jV�h�!:�*\3�Wǡ�fs��_\ً���Wb=�8�fC���՗����.�\��h�v��D�.��ّNn����g	�'ONkR�];����R�~��n�U[�!�uֺ�U9�ɢ�t/ң	MQf�S�>֯�F��Py�B�ٍ�ne�V����/s�i��0���n���h�-���4���/y����F^� 	"����'w�|�N�VcA�t�dq�+�ےh����L�! �q�Բ4�������6�t�r���"�X�!�.mr^jYz�VU�͙�O�,�=B�iO��T�o;�^a�B�l��:�ye���n6����Q�������E�܅jok� K"�cE���.��?�VQ>lִ�K�3�P�Ր������s\(�"
��OTk��ِWq:��f����Z�f�  ��g��Fi܋���W��=��&!_j�m�/�m=��;����z��\���Y/Lm��:[x�5~@��u�\l0�ؖ��Ow�>L�˱��W3&�k~�p��ܙ�
�1E"~btI�Q4�&]8ץ�phr�����]�PVU�-{E�Џ^/�ˀ�v��MJ߹K�$jvzg�Nh���zic���[��	�.�z�N)������j'�JHRQ���&���8������j�HF�ʃ،,ص�&���!UQ.�33QL�h��4����(�Ч�tQlB�m�5-/�B�R+LN�5U^;�'�����Q�zFk�������$)(�9l��<�v����"�G��r�f^���Z�vIM,�G,�d���T7��X���z�w*SV@�Z4۟1q)o�z�	���3�n'��D�����Ŝ��a9���҄�z���i���l�k������09��5$�O M�ZRkg�9�w��ܽ�C1^Ad�Ѣn�N�JaFR�K�~oX�.#[z���/qV�A��� #�q^�r�9%�������3���=';(�/�W�_�~2��8q��ax����*!y�u��@mw�0:E�PW��e��O-��)�h�\��Bn
 4j5�'��,q&��m�E� ��R���}�n� ���9�$KPfr���|��[�3=F�����Uv������T,(�S�t�	箋Ax��%��V�F��������N^�\��M4ֽ�[�.�}�v)���̰���3�L'���-���ٗ&�i�gi� D��36�X|�W�5���4[	輐��A'{�!d��dW������A�-�$&�\aS��X�vRX$� �ཡ��EHn���`.�;�
��7�{h�E����Ơ�u�è��|�V-g��
z��@�*̇�Jg�\զ�v8�B���Xt����ij�\r0�՚-��yO7T��s������F �s#����B �hA�e7�͍`
�u�U�zSosp��խ�H"�X�ݕ�Vp@gSv>8g�S��d��k\��_K��֎�9B�������p��"p�N}rՏ*l�$hɍ����!����BJ2۩�c�wrtp
��3��-���&��31S<YST���\*�����q>X�9���􈧳�pn�xgm�Tskt���/��k���-�벇�7��;�8Xߔ���mR�`H��X=<���6~�V��QT��U���-ُ�>VD2Д������4����v�� ���GB��B7����τw�Z'4o�>�4���("�;���Z���m�}�qj9{f3�+��bs���.t��ϫ�ƻ��:Z��,�u<n�⅒Uf�(��YH�U�+`m$M���6}�q��ȱ�>�'{�C�,#}�E�SCgg����'�w�H��q���x��wn�C�\�Ԯ��$�X�W�[��
�؝m�C=�v��N��?ܛ�V��o{���ez����,ڴ�IgQ]3^M�Ӆ�-��*M��71�:j�����"`�:gM�5�.�!��]��e-^F��j� c�kO�gS��O�3tƴZ�����}��v@;�	��"�w�݂�P=�‸��i �g� �6Gp#�Ч��2�W��OoP��q�^E9x���n���:�uWY����S�v������yG���Oa�)���W
Sv��c�*"���ٯ�>��@o�@��Q�i���C��[�],0s��'���a�ܮ�v�4[���j�9<D4�d�A�^=���3:k#@�0At1����e���o�O �Z�#0�XW%�!����}<h�/��*Δd<s�b����$��.��
i�g?�#�pA�Eb����h�M���u�+n\�F�@X>>���b�⚸��o>~���!����xM� Kv)����xHr�aM��(�a
�y~?-P����C����د�-�~,�:�`�R# ;F�zčR. Hd���T�~ �">�n�ULkE������c�X���&&����1ڟ��,><!zW�Ș�2)��"o��g�;� Gv���zU���ӎ��|�c����f{$��V2\ғg_�b��kO�.H@u5 �4 ��g܃Ղ��\��+xzn��bh�$_�w��FBe>� �ܖ�?j����
*�w�L�?CĿ$�n�1tޡ��2���!�����6�y�Hb�9���0��0CaE���6��-�OX��7����}ss8��h�� ޖ�k.��/^H�Cr1Z����I��D��VSQ��c�4s����;:('SH&�o�v��u]m����dU{g%+����Yii�}kyRў�3�4Y�n!�-�X��	�V�0śP�w�+ʒ§�k5`�|��o�2�f~)�?�.��e�_#mo\�K=��o��kz&K�ry���1��[�h�ljX[��U���81? Yœ$X��k��hG�q\M�et>�}Y�'���3�	n���*�ȟe�?%��":b�)���oX&{�||��H����{ ?����>���(��_�e�������#�:�@�T����S��l�~�ی�;�H�� ^�q�m������
GG�c�����%g/
CM.}!~���Ƭ��~��o��U� �q��71��b�N:�Aj�H&EO��:H�(�aUB-[O{ٶ�.�"�Hm��Z~2�^ �-�m���zQ_t��jޢKQ�
�����dYF/#�rfn�W�[�2U��aus_�_�0�c�y=�<��@hC���{=��d��u]�<�@�<��10fl�a��IJc���]MN2s ��9��"��=d#����ND��gX�g���[���l�p��m(s�6�F.>f��E�s��f76w�~�
������ЉI�w�2�\?Qd�5_�Fr��iu�A2��߉��2»������	j6E���_,�)�]94\#��<����0V�x:��X�k�I�Y8Ot��?�=�e���6~K��#hI�b�E(�������䋚�r�m���}��%?��ɿ0�J�9'%Y��1T�q���ۺalL��o� G[��@�N{�3�Мi�OS�~���jk J�i���UR���Z��ٗ{�)xׯ�v��<V"����+�� ,ƒ��"�6�˥d&��?D�2}����P����`�Y�rX��,������x���(�Sy!pQ�ɜEv�{}	-����U��txId����.^$���Q?�t{=�;p�������O���b+t^�~���S�\���e��N�(�"3�t��pԆX#�Nx�}ťw���b�}b�C=bz��@H 1Gñv����@�a+j��w��K����zM��(#8������\'�5P'!�� �X�I/�\�㋐Js�Z�dL�]T���:��Ur��;�[%��p�혐N/�?-x��� E&�������|���MS���O�9�S�r�=��᭴5//v�}���*�R�K�����ʷ��viO
�&��g�����5LQ$���L���=cڛI�c���v=�a��ߗ����*��G��w����F�����'&>��&��u̔7xv���bmbTڞ���ȏS��'l3j�.w���?�6[�V��|�p����zgJ���d��T�����p3��{B��ٓ�0�G|MXp,��̀҄d��WF�.��	�m��L�D9�yW�ǒoG���o���xL�L/b@d��Ə���T��|��p��pC�$Ã�A��W)�90��d���&
�pj9�Q��h� �|�4}��K�-�a���!(RV೶�a���Ϣ�j�Ʒ�L�a"���i�%A�H�&�3�aݸ�~$JJ�G����_���Ԧ�T(Nۋ_��7�e�!��|�Yl������r��+M��ߝ��.�2���<�2k�'�_�&s�I!g�#��������go�+Ct��� ��3[ N"�DK��Zs�N:�.�鴒����M�H6�o�A qT.���ݴ�3���$�hwL�Qre����
�vἕ�ѯy����1fN��a�U^wP>�	j>�H�rI��+0%���v���_fG��bԉ�A��P���bY1{�3џ�:�S����]6�jy��1ҧ�.���77�5����ċΕ��Ux����	��5���E\0䫥S�����b`�����7Ѯ���3�eٱ6�w:.�8��0S��|���מ����KN#7�咰o{>�LU�7�7_�����E����9�3z�lp�B�g��?���zp�2�Mfjc4~B���ͯ�[�$�4��6�_\9�_����������sZ/ʗ�$�%��6���������Jm���Sʓ��~P$*鉽rOX���ty��CE�1�-�.����@<`׏,'�`*�VQ��U�8=�}�fˑ-��VT�_�%����t�n�Ak5��$�$��U#5k7Q���"ll�`'ӏ� �6O�ӶУ��Ab���j,T0��v�)1�C�t�i�G��܇��!+-H3df8�F,K����]����,	E<e�
��_���?��e�F� st�����EP���+��+�G�!T7�>�(�ܽ?Z,�����o�	�ᕦ��Q��ȓW�u'Ԉ�+�������bܠL;�����t-Py�1|��4�Bh�[�T�>¦����$�Rt!"&5����'#��PB2"+t����:��Yף��"`1[:D��D+^�Zƿ/��a(�?�I����@���ǹ�~k��4iB=&����K���	(�Wh�c'���|�vi�co�)%��Qђ����B�6^����yT+�ĩS�r2>�^��G�����T�r��eR��{`ğ����u~�a�&�pf�4����`UƓ6pZ���N,H�b���\�c&赺�N&���1�?���l4]�}К �b�P�{X�#��<t���uŗ�(�g���C�����ޙ���s�{WPt���n�9*���`e�#c,�w~pB�΃��G �^��h?>*�)]��@��|��	7��Z&�A5%�z*b���|>
��LXo.>Տ�� qY�T��a�^��.=`��P݂�e�ë��zހ3�h�F�;���	����uj�&��s�D�P�!ƿ����-m�3����>�ސ��KÆ�h��]����.�S*����3T.z�#|Ƈ��0��m��+iƾU#��������ت#���4E�b3�Rx1xo܍H1��
8eI�J�O���K�UfC��eo�Fe�m�J��V�W5pr��s����ތL��M(��s�X�Zی�~٘����<���&�<������}��EL24T>����F���|��4W��.���c��Ɇ#��v���;�%+�_�lu1�̤��#R�8P
�!�X��M�۪�&D]����h�Ÿ���!`V���oC�=��ܙ3�i���aEuak+<,j��Qx�q��H����d�RSش���
{C[i�'�UV���+�-CGN�32c��h�;�ˮ���)2�G�g��}�������0*�}�cD9��B��k����x���}�������ݔ��5ƨ�q�X��B��� y�����B�7W�����bL��#`@�o�c�0����B�<�L�;��+5�	��&bV��h'�6WQ"%(X�Ɂ�k���gL��|`�� �-��}�y��=}��b�\�X���}���߿������C	C�!���rtw�W�r��P&��%A���RX�E#�:��9�m�D�2���VT��Y�W�'D�ΌׄW><6��8��|�\h$AY�FH�������2vrAvlf
Ԛ��T�u(WG# ��%���IV�`%v�a�>��%��;�`��3�M��@�@}���g�K����Ey݇k����Qg�_�`ұe�1Sv�y�����f��d��,��	:U.�j��y��<p�7����a�g�(s��D�&gT���p��)C3�R�A�6=S&j����f��F$8X��1\t.��d<'#檳�j��M�=�YK�V2P�9
G�IMQ��I&�'"��p�q��F�;IW�?9%�k��}�I �O��������^)ٟ�A��V̒��⿕9a���5��>�mqP4���Z���� ��{��,:T�kxL�,��犞���&]l�R��?��k�`���%�8��QK�˪(H��*�?F<�ѣې���%v�o���?�]'o}���>V#<��.�ǜ�[!��� �/�
�gӫ$��Z?#�����p�/n&���-�ȖA��W\1�-1�[�A81�(��m�Hw�}�K���e8)�%�1��Z̹��"VB,�[��B��4��,Ͻ�<,߃;�d�I�58i<�q�j�Q$Y�,��zF������]�`�'�$Č����u��ӛ�,ⵕl�4��BCB-�W}�-A���U�S�o��Î=>etQ�@���(Ǩ����<�d�`���\k���jݜ-���e�:�4�ui}���J�|���$8\� 56�.r�rK��q�ﾲItԣ�0����B���N������	�%1�J�D��Aa��ЀM-E�r(v�e*�u�U�q���C��+\���؊��'�5U���n��� Nt�
ǥ�"��)��S������U_�C�!�{Gx��a�sc�3�I@���N+�}�]�;qd�R��1�&���	ʛ��~5��kb�M�r�
B.B���2Ґ%M��.|�*r��������C�t?q�KQs"m�!���%����YϺ=�@L��.d}�2�`�S�|1���c��6t�m�D&��s߇���Ff��2牡V5�C��s�P���uz�Op}�!�����-!G��8~� ��\P4��v����3?=��V�[�|x*o-��9��%������MB�;�.�#���_L�gν�3�)*O�.l�`����mk!����8B�t+�l����v�rD�	Za�e�]���텓ۗt#��+���Y�@�XB�w�P����$��p,1��ZE��n��О�Eljl��Y�����>Aٹ�&~��I�tXm���?'k=�[����Τ���$��)~�N��RgSN�7����sOm2^��[p��F�������"
6���\�T�yw�e^�⩹6�.C!K��Tt9��޲\�A�Zת�����ڍ�H��Ѡ���a���/=��$�ot�L�`�s��k�G�� �2N\<�0��Y�+/��iWw4d�q������[��q�/�kS���+Ay��=O�+>>��� ��=�,Z+n̪7P��}���P�UsKz�G��(�*P��
өF�.���U��Nk�M~Q�����?�ʌ��7��*1����af���� �r��Ml`e?DtA���~}���<�)H��V|�-3ޤ��V�4'��vk�*�����cWw@M���� ���(r~2f��gn�_��Z�fPi=�f���R��U�.���ꀦ���F��*���g��UQ��;^�pI���-�:�Q�]�_�ڈ�&/�ѓ�\�3%�չb�� �{�Y��4�4l��/I��R��ο/��y�l�9��tn'F�r����:%���?�*u��NW��*L�50_�1�(�G\����]FzuN�$��Cn!�f���d�@j�ؒ�lI�\�E6�	'�c'lSP>w̄�)��f2�OO}�`i[C<ĤM"P|ٝYC����Ec�+H���V���R�.R,���l
.�w��m�Gr��*�(^���B:��ܶ�"@ �s�F�)7��Y �2@�gL��){{�r1�믙�<o|�n�.b��uh�5���:Me�ϓGwu�Q�ay㜡b�3���=H�,�H�r���ʌB��x�b�ґ��=uGT{�
7-��q����^A%3_�
>�W&_��!  Q.S��$3���IG�D�<�� �8~����E��<6sY�;P���R��U?���*B�H�N�,�D+��b�~sN�ͺ�AO�1�/�� a�k`z�� ����$lK�[��YyW,:^���/�B#1�~,�'L��G��Ό��=Bb¥��j������"/T#W`��zlF��0��ɢB�G�e:z���b֣������g�j�Aa..�b�7yc.ʺ�E����߁���Y����fbBY*�b�:�l���g��� �����M<(W�;��׆�;{U��3l���,7��b�ߘ�	Zd���ȝ�ȕ=n�M��5d��9�0���SD�剥���쑲��x	i����\�0֫8�@��g}��O;P������'�Q��"`!Z%����+8^1�6mRx��?����NA�w޿���^��\�݋�����Y^E��>�[mn�"�`�n�#_��{���)��¶v+���)�\,]v��6�|Y��p����Va��Ag��B�0�.�@�0�ł*��ru?�'��b?�t��Ǣ�����)3bU|�L�{������ ����i��`˟��I��g�zɇ}6�݉-���ř�z@�Hv'<Eh����@c��7�j�ɾ��:R.Z��d��)��!���v�^�_�v)����X����&d��qy���������ـ%{ك&E��4\���T�p')iй�s�Н",����M���K���׹���[��C��Y7=�m%������E��<��d��z֦����ޤ�{��<�ݶ@W����A��p3&�D	a�`�1�Z�#���Ìu6�e|��bJ���.�t��;N+�BNm�D���6��eA7M=�6_��~���6�������U�OՂ�֑������n�����׮c����{[�X�3��\5���0���""�����e���?���ɔg�y]7̀�Ϳ]���­�HJ�P)~cѐ6���ǔ���eu&�B)��E�:��fTOh\tU{��]+��5�٦���� �*�,������ׇϔ/��N�M�Ӽivf|�=iΓ^{����^�����������E��N���C��APL�h7¤�����=C^�l�)M��sKv��v'�������E�7%a%WB���F z�h!������[pÎ_w��>������F�z�ܻ���eFw1�L(������CD<���?��:a`���Wl�Z
OFrӔ�.���;���<���,Y�
�Cb{;�tdZ�ߊ�ŗ���c��}��?���t�]]r/0Ȓ�ta�q�3Pլo��F���_�\�`�ȫ�͢!�}a����u��&,���\(µy�
�
�F�y^x���?����YN��oҭ�K:�� ����Vl"��8���'I!m��p��h^&sUz,	��3�N��>�@�M�(�Bjz��=����d�m�*Li�Ƹ@�3`���\����z�N��"+Ms5�4���ω�����P�]>~��y�"B�:dY��c�������:�7Ôs%�� �����"ҿ8�s��m�׭�P�������?�s���H�ofU�3�WYN_�݊ �!���$C30vU�bp�M��,��XȾ=����._a������h����?����h���R2���8�)6��T ά��H�}����"ZQ�|��l��yJo��Rb�d����F�S�XA�n�����g<�݅���62 �����n��5�x���6M�m�ewGiә���_�՛L*=�2�nGW�$S�D���r��P
��5�l��1��ۘ���q�y�:7�6^���;��?36�9�MɔWˇqG�2"xT=�;�*ҕ�+���=Lw��N�o����]�4H���Y�Y�/Ĵ��"�4b"ӺN��̛ P93�C���4�0�.]�s&��?�Oƈ����z(������ל�P�i��V��&T���G��7�b]�:��`�˭^���X������%�`�8}1ϋ��l��C'��Y;�gH�:�P����09��?��l�P(.�o�%/����gP��D����n�	�����Ҋ��4i]Wn��]�C��sK(��9鱋\7���N^��@|�(}�Iq���)Y�5�[����.9�f�M�U��Q|8��@���d�I]����h)��Y��a����{7I)���W��|r�3��:��Y�%��8��O����Ud�s�D����z3Bt޼���{UN]���gkx�g&)I�L]�gw�������=��5���|C�K�����Y��Z^����bj.��r�{����X!Hji?��� CC�������<~z3���	{R��>.Ф�6/k�mw$d�|Rŋ ��G�w۫�5F��kJ&ҥ��Z��4�|�ip*>�p��O��u��^�vMCpc���o(<	G��o���[�d�[����)�[(@�4���q����2Ƣ�g� �<����$�1E�e���B�/�&�/��(����v����B%��-^m$�m4j
�����Fk:{�]���s���/3|��L[��
&XQƪ!f��Õܸ�gq7�B14��DВ�S)+N������4z��SEP~��S�wu�4�|�����j�س]-�Y���, 3�;�H�Ϟ��JL��y�Y��_>��]�G߬�c?FA�\��S�*��� �uU̽J���a_���^V�[�F���Q�s������7zФ"���:�.�!j�� ��i�:���p\0#6��9)�Mo'�e��=g�{{�>��rN!�WA���2�h0R=׶'.܀K���^�ސiq"f��S����tcנ���g͒�#/_7�e�u��Ȃ��G�����0BCC�!�E$ީ.�Є$���#_��0����Y��y��~fs���B�joƭ%��B��۴[�2k���/,ڱs�V��zHK�$�ap��OD�����I?� d�^a� �a�k�UV��w�k�I�
�����4h�$�F�<��R䙾�
��/��o�.u��k"%�����-��V�v�����
��9֦U旽�$��,I�Rf�\�D��f����%b3Ĳ�Bn0`i|��ݥ:�J7с:��c �@|��NJ��C����z\��l��X���C�YN�,p�J���*���� i�>)A�8僚f��ǰُ�H��%�e�߾��آ�޻�#pA�*���1���5E3B��ǽ��=�v����m'��4$�y9Ѱr��/���cZ�f�3ЗGc́:�T�����e���[���b{�y'���1S���M�o�����t��<|f�Ep�Y������,V���#L����aTq���R��K�m����2I��{���������6���X�=�՞>Z}:R���[�B��ۉ�&���axWP-�d����J�K^�ހc��nCB�+^N~�+�^B%B゘�c�9������j^=�ΔFzYg�����]���f�3K�.L��$�)�����8�q�<x�n�9�2Wʓ>��*��%�
_8�)r��|�2.T�<��LZռ�~be'o�|�kʓ��|ⷉ^[�1m}�� �l��.�fg�>k�WV�L�1|�tM��ٰ�g�&�
��9-?7�A�%W-* <�̐���o�4�ߵ�Wʛ�De
�=L5���P�[����7u�5Ἧ�JQ�ف�8#J�#Ɏ�J�ߒ�劣���"���ԡ}y�hDc�<nr֮��NwG]w��H� �{�O;���&�P��И���J���� �\�.�����J�o��������Ŗ��IJ�YĢt��!�	'JEĹ�qJ���/����T���Uσb Ӳ�����v�v~��t�-��6��y���`����Ӊꡑ*N<yJF`gp�g9ʦǅ������t��,��{��x���
:J��%d}�&�'�V\��("�uu���n��j��h�t&�&�2k�j$EB�ry��ULQ.L����$�e�So>��O�C�=��58o�W'r�
�p���Vht\'�����S#�����Lc sb�����o1��w��wT��C��i�f0��"L��D��V}�8�& ہ}�wщ�p����ۻ�эay�x�CmiS�t@G���Q;-4�Ipٷ0(����Jyg�^Md�
!�W��5���S���e3Vt��Қ�t`����<�״�ˢ��A��t�x�g����_�&|r�<��Od��9��q���U���Nn���hHh���?6qr'7�+��p\�A�dv�sh?A�M	0�d�1~��IUO���Q'�ɜ*������
_���j��`���w�r{*T ��+�/�������U���;�Q+>W�pG?����֘c���wHމ�\Y�º�ՔZd�9��a���gӨ������V
���:�͉�o�e��ߡ���/����o�l2�U{/��](��R�t�A#@�`M��e��ߺ������t�ךFo������J#ۗ���G�wWm�
|���+3���e��1q�y,=tL?��y.����Z��AP�]g�_��:���~[dDSꬻn7c�Gŷ{�sR����`SMK���O/�:���L�\0�����i�K�u���uvS#�G�D*J`ֶ�|�m��o<$�A.�Xw���q#�K�鴥���`�F�Z�p^����vB���<�-�8%O���6{���+�O������N"��zV�Fm��dC��J�sǷ��_��E�K× �O���|�Y�K�ճ'�:ĕ�Q
��ˋI$��V�M��i���O6�]�&#��.4[�Z	�-���nfn�*ĸ�`�b��3۠��:�R��v٦��V��|������x�E���g�3�Hb+o��u�h�C+H�20��c>��,[h����7s߽t"����Ճ����Q�ֶ�������\Ь�ݞEd5�@P��m�y�$C��[�cy�f��Y��d��M�ľ���Т��� �=��2Ǡi�jmI�X�7��-����sH��,I(5��R�5'����e]�*1͙����yt��-6��i�ya����#S�3T��ܦs1��v���Z���h'4R[*Y���Fw(�	ҕ�U�Y�	���iz���}; �%�v5}�8[иO�؀R|e�k�?3��Εر=���U�HL�븎�y�V�[�G1Nnk����S^S�)�7��.<fջ�4�BBB@��񟗰˅�}�7�8�r��� �ȅ��I	����i���s]�'Ot~��^o�4��cZ\�H�[�ݠa���ZN����O.M��kV�7�����SLS�o����6�@=��hU�����~<������\�gL]��&��03j|K����x����)U���]j���E����X��*��������X������J�a/`�G=u�d"�b��~	P{c$�#��������)VU��%����U���Tg�9��Q|�e�29��ژ���0O[�|Ʈyy�&=�%�jۣ��e^p��ţ~3��5刣?����!DM�)U�gTgEy	Q��~=��#y�Ֆ�@"_67�`���?���<��w;˲�e�)!��eޣ�ef�'b����]������:T�{��B��ퟱ�Y)�k�ߜjq�_B(��nJW�<ogW)"�S|~�<H�^�c#۔7��?�8�9�U�`*u,�-��r��8l�V�I sݜYb�g���6�1��A8�rȍq��0��r�r��z�?��G�⠻d>���w0������@{_F��Xg��V�x������,�A
m����w���5>�義�k�Nטtŭ/1Ԗ
�`1��0٨�!LZ{��N	�b-��DP=D�[��H����؆�/��}�J��P��a��䜺��ZJ������7�|��#�L����n�5¥�.�}_^�S>��e�]�,*!۴@��ߦ�]r�vP�\��w�U^����*�WX��h�"��=-�d��c�g�G��f-x�9
���i�
~��EGwA������O���	�ֺrz���^U��J؏:*���9�g8h��Q��_W$O�V-;�ηX$IK;�bG	H'}���Jm�¢�^3?n�����G+�� �d�6��FA;K)��w�u�Rpc�v��O9��e�E�H�-Ft��o��BQә�bn��U	�,b�PL"��`�*\uFͅI�+�,S����\������~�偰�O�00գ��_)�لo���݊t��/��u��̺B�z�u��e��c����6�����(w|ĕ���/����Ơ��*X G
���)t�hk��?���$Snj�%�����O�I�{� F߰�u1EF�L��dm�-���{�kH��I����5)
D�Ǿ���]�U�N��l���C��F��K�w��2TR���#&B)�TІG{ѐg�g�N�r�?�Y��N���6!�h/0�LZ�,�q󅟸��F��u�;����Kv-@�J��M��q��5��]*��c-7IdǮdZ����\�ЦxI5�,f	O�E�/�aIQ��Ic��}!��ރ�ꇡLp �ǥ�s&B�\���ʛٰ�����y��Ѝ!8{�ܛ�ztC�������@@y�d��4D����F����u���xQ�F�:�wW$�`/,��W��M��nƔb{a�;��l$]�M��4�����H$����x��&{�|1%GuE�F$�]��:��o,T�_;&�ڬ�,�N�T����y	�]2QvƂ���c	"",؄#t6Uw/4�N~��U�-��f�#o��HR�r& �ܝ�GA���!AL��E�$��>��$�%xhX���n�zJD_�^�����	�;C����N>X�E�M��pL��%�=�I�*��Lͭ�@���dm�&1p�R!�1���Euy�2�0z	,�
5v�%�'M�l*�gǝ�m��!��`���"�n5ϭ´�,/��b��	�7&���Q7;u�D�-��n:͍�Fo�<���k��tZҗ�������7x
��ύ,�g<���x��Yimj��.vp���Ea��STm?$>q�µ�.<[d�nn��y�v���`�Ǣ���Q���
��h�Ȟ���K�|����*a��
�� ����s�|�-�繌G�g��AY�
��^��"�V��Jj����vso�H�,s����=��%7���C���N��"�d�QlP\媋��`Y��h]�2.]�^i�v~�G"�^�6 zq�T�H��G�U��h���K"t_LI/���x��v����WSI�b��:&�2P��D�l���3���m�p�IՍH�ǪW#������e(v m������!�X���P��1��~�$���c��:ma$ńt��""�黸>�5|���EY�/�BHY�Lv˼ŝy�L'��4dCmg��շ��X!w)&A�����rit��L�8�-���n��J���OH�o	�v#�1{�kɪ�]�d�o�'�{�A�͵���m�vf�FY�h�a���*+�bJ�`e'3�,����F�'W��l�Mo����ɶ7X{�v�JGyF���x�]��τMMF����z�g۷N�wz���u&C�K)�!��t��&�?Qd@��|��YF�+�Q*0��8�N�hO�R���6�y=h�"��u�Fa��;�2:G���(��n�ا�]~tƺ-��bU� �@���؟Lʊ�5��ܴ�����'�	�7JHg}�.,#��M�/���XY� k�a���C�Sp��qP�Pav�ݠ������*��3�u�au���(���ΰT�����r;=���S'��3S��r�qu(��5W<�eD*����4`~@NNZ��8+58S+3�� �l_�	�w4A�W�1.��t�b=����C+ )6�$�Ii�����|}D��H�w��������(�:��;E����ΪI�[�)�k�ӝS�;;p����k����'����,T|����ֽ��1D�Xå��:�5^����� �Ļ~�D%貭T���*7	��)3��Q[�޻G\�~�m���jQ,J����nj�-�X�6*��K���F�v�v�d��4�e�s�#>�Z�+�����*�5H��h_���=@Ԍy��B2Ȯ64H(����S1�2V�C�V�bw��W�=qL?���5�K�m.A9�3�<�Tw���r7��xr�Z�,]Oy ����~�T����a��ە��Y�N��EK?Uk9c�!8�B��\�b%32��������.s|zw�g)��>�fE��|���!�=缞�Q��aH�@Qf��d���JQt=O�'	8�̺��:U�b�1���U"��_ Z�ޜ����է�~��0q��2=�\����e%`\�d��:��v�F���T;~'�'�h*q�m��!�|7i��]ϳ�?sD��}p�v%0U��l7E]��1�BK���$�<��0��R�LM�~2T��~	�bSdD��M�;���H�+�W����-`m��v¹߃Dn x�j��c���|x��MK�d`��cS����כ>� ���Ġ���q0��p��.���2�o_J]e0ZӀȾe���g'$�0�Z��;ń]5��݄��g~S�M��®ҺkV�&x�PK5��rKr_�d�>�-Й��~U���W>���7,�n�k���I]E�'8g����Ǆ�BI���[dx����i�/��D��A�f�� ��A��uOM�*��S��U~� �@�$e�Fjj{��T$Ƭ��;-��S{H�HpNϚS�Z�	�<�M�7SNW��s�LȖ�ϳ��wN}�|ĉ��7�84�2�SI5���i1��?�s���p�#�U��A8�P-�ip��1c�ˀc�CL�=��<�p,�dr�%����	6��;�>FL�ً����&my�~5�2{�Z��sCq��+�5Pd5��W=��HIU���-�ԅvWË�^
dǂ63��56�*��F�����D���`��� B�b�cL�������H��)R����ފȯ���S��W? v-�c��ȿ�2"[�G�:�Wwg)F��#�W.B��kӰ5e>{��up^�.��v����5���E�x���Ҝ3�,�`����cn��2�"4�BfV���#�0��S�����Wj�0\�Q.�~�vb�]U���b�T�{�iw�~����� �XU��rl�:Z�&�[2�Х��o���5��6��j撠�;}� �g�q� �'�F�K+ιt�0(��cXm˾�W�J�X����.����27;b��&�j%CF��C�њ�nZ���`DLjJ!e*_�K���n4:#;G��>����81���]U���SI�e����/�����^+�4'o���G@q����52cw���9f��r�����ʐ�kE��ۻm]j\����@��s��GX�%�[sF�L\�ܸ�#�_
���Q�?��c[��� �2���4Ţa�A�<-�l5�� �#ͦ4-$W���`�M�N���*}�QLk�^"㕒��C��^Ȕ�z� �KR���.�z 1�pH��;WR�퉪�/"��B�.�,1��M6�_cu�3ɛ����J��7�TҞ6=O]����"��Xځ��Ky{��v�Bi�2��M<
��T��4_���p69�G��$Z�ʷ��~׿���%rF��\�t���P��O�1�A7�#FԷϘ�
���J����;rA�%K��1\H�~ӎ�`o9�S�jH+t���:j7�\'+#�r�˪L���^���0obہ$���y�;$^�B�5S2���==Ԫ��I��f�K���<����e�|IƠvB"ꤐ��U墖�fX��'F����Δu_ c�	��Gb��HV8��eIfx���~�:owh�W�T������l���W�u`�l�L�4�^�NtD)y*���:��Y4��
�T���i��cB�w������b�ҝ��R���-I��d+2(}�諐*X.�B�j7������`/w(�3��97"{5�?�ڻbR.�g�aA��|X��e;�����-;�\i��b�ٺXP�cY0�K"���oBG�!@F[���T�;94{ ���j�F~!e3�70����o?U?j�x�8�ZD�팴�w+0ӆ+�����
��{'r/�f��`p����δ�΋�'Z8FF����~Y��(�w�G�i���"ݬ�����0�)��@��)��������0�f�+�y����{���S�3�i!U��N@�">r���9����fS���*�z���Ag���B�I�b�ie��ڕ� �sP5��&���I�`������</�0Ս}�lzx]脺g���{�ō?ۄ(��z��tk��!6Va��lyg��뙉�B��k�Q��,���i�Hq�\4�!���9V�6�OuS���$�Nd����[;��d��l09��x��n*�|k�p�l�U���twJ"�\g:l	�#��̈́�K��ƿ�7��U�8���E�W��!�S6�x�Aө�2w��q�$q�+��c�m=d�vz��y��]���n�.�"���ۀxLE�@��:�1O~�Fұ��g��η�T��h?'���`V��<,�dD0���[�0-�R*l�z}��!����%�"��v��4\Z!$���w��^����7	cy�J@�T�[x��N}�#V)1��Ѓ?U_�v��j������߅?j��B/\	�;���kT�W� CG�ͅ�VU�U�T�wA����h�I�����T�:W��CoR(���?�'B��:#�9���Ka��%h9�#J���� �HHє��|x�=o�܂ע����F�N��Qw�hO=��7�Ɍ�f=�䶽�3��7��`=⛀cLg�jQ����E��[lR�#�G�Q]4VyB��5B��~��9�n�Ů�u�A�g���A�1W�P4�hh�;���;�v�$�X�乯�I -y5q�ؘ��s��9�u��L���pS�]J'RY+�Z�ҌJM��Z�v@�I�����7�d��7��c��_7CO,N�a�#8��Ѕ�3�d�׎�L����1�aj~:�g���ѐ��8FL�a�/"� �G��ɎR��rGΌ�Go�SJ��b��s�>����G��P�)�?�,:���>�	��&�������f&���1*oD�������'�C�����Jb^Y�ɻwdEl:q��rgz��ͳ�)�7��7Y�7�� s�ܱ���ޜ��M� �q�tnO�ӆψ�S#��l9��jp�Vj��S'x��G�}Y�e�$bh��������"��mz�(�H�Q��i�-��i��k3�1N��g��R�x��y�p���T�a {9���t_��d�zg�2�P��;q�]� X�'D_}}�lq�7�%ͼ^�z=�k�Â�z�<i�Pߓ�s�[��RHyM�~�������O�F핵�J�����E��;����).�R��RODe;�RϢ��u!�=�I��V�33����򌝗�D0�{ձs�|��q\y���?�-�o��%a���]�T�ׂ��i�tl�~:ד��dgo��Қ� G�\��� �?�
���Lx'�w�M7!��ag��?�jS�6\�h��B��FD.���uQGA�a��<�h�]˻N�8����c�v���]p��_.� j@Z�jtڂ�W>��5�tİ{Ti���{�op�����2���ӥ�a���:b:��c��F�9#im���0Z8�e��9�J1��}��".�FJ[������K06�p��M�kJ?�b]�)@g��>Cx��m%~�G�s�%�Ӗ�Ҿt���-�>DI�MB��%����:5K��=�� ����>��ԁ����>Gu��2�SI���#9�&i����54Ñ���ޮ�a�����~66V��C�i۬�ic��Ĕ�÷���*���p+W�Ƶ�r&�4/V����P�>�{p�E�-EK���.���K���Ȗ�<�V��Z�	���%���u8�Fݣ�R�~���U1�~��[��my��ܒ�h��(1�y�H����S��١w�6�̆���Oo���Y�Ѹ?�&c�����y�-�<�h��	͑���{\Q`��z�-l[NU@|��Uי�� �H�j�����8{�_��GuDY*����_��s� �_c;�fE��hkI��rQ����ݺ�z�k� �@R�E$i�jQ�vlM]��j\)&�8t��i*F���ڀW���'"�uu�J��]�{�3�c��TY@:!/p�Տ�OgE�-ܥ�VO�N�Q֧�)�8�4�?
����Uzc�W�a���<�>!�]n����2�mԺ�-sL�ʆ��%�\�`V��Ęl��k��0�� ����,����g<�����l �&��a`�n��Z�q��-Xe�&��#���9����~��X���,�\s�?n��ڠ�9?��Cc#�r���,�:�q�v'�/���z:�BM�z�H4�"�z�̣4������;
>rL��S
�W.��څ��<; �=2ޓ�#��q�װ�F,P�4�d�������n�`�P�A���	��_���o���>�2�?��"�>�V	C*��"��kl�4����+51�OU}v�[��#�`T1P�����!�1U�h<���C�plZ7#��������e��U�1�j�fmF֟�o���A���~ �Pa-�e�:��q�R���o{�m��BJ{/��`H�=%1�ct>��Y��#ҋ8b(�r���S�v޽}����P��x<c��9��� i�`˭�H��RRK��%\��u���s-}UP�Lȯz�L>[Y"�ה# f���=ċp���*��')��k�$"%�T�Pm�K8�`˫���ɵP!��v�u:	z�F��5�f�}�ve�o�$A�+9�QZX�$��ј��!t."Ӫ���j</m��U����C��;��8�eK9s�E������B�E�3�Z��+�G������Z��}\x�%��Ʌ��2��S![,'+rm�V�\�����6��=�b~�����;~���m��q���K+{�B�Kg��x�������w5�z� �en�����s�	����@��\Jӯ�'��3P���9v�cf �I5כ�!~��J�8.L�ޛ�0.M�i�4�,l��Y�i	�ȯ)lK0� o�"��=T�)�7�LX����W����fVE�t��T��[�S1�y�V&�
��sq�t�p�X�-1ו����Ub09��5�hr|�Th�j��@��؛~��u���1���H8�'�m��^W��F�u���9�x� �7A�6�tzz�`n�k��\� ���8,��z���¶��T[�Ǟ��@����o)���e�
9+1�f�o�}�1�v�s�ԴQq�!� Q��Qm ���
"��d�/@�b
J�6#O�S%u�7�T7@鞝�z�������|'�ȳ�� �� �+�m��Tf�m��h_�AG�����0+y9�����^7��SxQ����|�z���D��X#�jM�/�W1�|�2'�������~�~+�������-p���Ft!�&��vf4n����<�Z03]x�p�r�%B�(���� S���Ǭ��ؽ)ъ=���.d��4��2_���<��M�|\�i�`�V����\zRl�*�&��+��o1�� �y��w?���b�R��(�R��5����l����2�E9�u��RD@��Y�3�O��aߗ縥'��IGq�$����s�a�b��P�lIv-<�67[R�W���F���Ԭ�ټ���K;��y��!�"�w��c#�#4[Ùudxɶ6��O���j�^���#Mo!� �]d+i*J��?�0J�c0�	W`�\���%h�]ʑף�� ���-P�����?�FG�pL��)����a��5θC/#��8F l0����V'ɾ(��j��}�{����;�*�'�&C��{��ȕ.~f��[�aD�&�Y�!� �tr�R�e}��p,��S��=$�A}�H�]�A�6�ŎZ ���'Զ��֝��(�XC9�[!� C諬t)��ouі/�.7.ZLU-Pm��7ڛ�J\�Tv�?}򦺱��F�d�����Mg��Q��+"cO����	�Az 6�u��s�<���7y��ŖR�l�5��V�l�HG���B{����:��S&��� pt8e?D�v�x�K�Ӎu� uA�~�%YNؒ/DT�i\��S0G����.�D+�^nKN�֙RYYi��]�6
v���w�?�����x��}�	W�/Gv��6(_���Z��h�~czw(K��D��=`�_�C0�}����?��%y��e���fN~BG��H�p���4�QN�_�G,� �9�2��	I�1���J�31 r�h�*�xpn�+�d�G�=���y���?	�	��4�V=+��uw�Ś{Ʃ�Ty�B0�i=/�4�U~/8�,|����.o�|�)�7+����A+ĖG��	��%�U���PeH��V�.,�#j�!rԪD��`�&X,��aP���j�g_9��?�ึ��?pY҉�RFl����Ӕl�L,�P��;l%&�`�#���b��q������������yA9�F8�6ё[nÇ��!Z�����b�����Splg�~I�D@#|n����V�k��~��D��K�v�yK���V&~��:��$j9��Q�U��Ԋ�.���|�z1�,�:ׂ����`0����TI2(�p� 9��[��	���sO����6*R�w�YS��\��eA�6%�\�y�/]�Й J��7����:U.)�Z��75�3��7��p�NJ��$��l�-��}%���A�^�G�l��Zy~�8I�ƅ`Fd��l}`�J=D	W��x�����J�&�]��F�hЊ�󁣫J�Y�.&ċ�4J] v�C�(a���ͩ�kj �A��L��+��+}��n,{M�)Hv�����W	�yf.��H��~�M��J��D��g��r�nT�����Hg�VP�=6b�,��?<9�XeƝ�Y�SH�Y����T4��J/@�9�ai��-�r�ǿ_P
+��ԳI�ݜO��w��;©�}��Ȃ]c#�� ����%��c	��4�Y��/�癛��'���X�mCo�⃲�R�V�IO�0��Pc���H<��g�Mx��`b�{[Gh�£�.���*7�P���gj���|U��{�e�K:��ם�A�e��m�PcФ���%.4�
�nJc|x��wI)�w�c��b~69R�h/(�2X|BsS��H7+:�o�f��n��p��W�?�j��Z�@�k�|04H���~(<�'Po*T�|�3G@���L���+P�}�a ��m[�m�Nȥ^i��2���2$�=��������]0QgǷw3�Xk>7B�D��L�!�v��㳬t>�Ģ$7,�m����p�)��A�˱��h���z9�t�W�^жf�B�ԛ�R�� �})'i%-�գD���|z�!~:�F$z�]��h*��J�M�])�置'�y��OH���Y��HtMK������$���S<%�n�N��ڡ5S*3Ô����YMɡ)���O�s�GK�1$��5�����M�W���ŝ���XH�LNkQ���E�2Z
4���V~��1D�����>S?Z�u����ǇL�;��u���z��^�`9NRrY��?tz!u&yy$��/�7���cMk�4{s���#�u!I��h ���ӫ2��m�4`v0�Ná�u�F����'�KԮTp����D���s���N#��7�'�\T�@u+\A���EI���v�y�ʏUc��2�u�2��B��]kqHl&ն��-٦Y��?�Ê���p�
��k�;�j+�#�b}�s���l�����:b�{�`�-w��l\�)�ʀYN'���毚���nB�zO�{\$�~\����&�B^�v��)"�{:���TzP�r��C�(���#6'�\��Bs�����Ƒf���X�OS>�ڢhЛh��	�S�h��Z`i]n���60��wS�� >ۓC�V�T3_pH|��&�:sQVB� �q���,_��n�89Q� gl��=�$�9����2!�(��l} z��,��'Yni�T�Tv�_��/܂[N���M���W�N�	�fΗ?��ra��Jc_�e�J����1,�TH��,z;<�<�[�	YD+���)C}�S�0�yW�4���tx�В�8ר�' .9Q$>Z�O0��޶(�q)с��l1���1K��A����P���iP�l�scћQ �l��������h�{�A}Ϸ�P/~'i2D��B苅�uB�Q��y�s�LZ����,���ف��2豢�s��Hύf��ny �(	��@_��~ 0�g����E�y�c@t"���DL䗛}��TP#��w��l��-El.l�����$6� �T�%
��Kud�����T���Ȏ�r������"4G��|R&����S�f���#͝|����<�Z�1���Al��:m6�u�D&����� ��0����Q�Ͻ����y���\n������.WU�������ͬ�f[	υ�ȓ�}�t��;;p��?%��ƁN)_��H�`E�>�y>���QF���{����{�YƼ�{�熄%�5|^Ȕ6lb�`��BN>KЂ�=+�
��95Ս����JL���������g�n�cV����~Z���4��D�(��)0��-f�%Oc�Pk�o�w���d}20熨K��T I�ف�� �a��-�@�Su�6�I)�hԏ�~/��"����o��Y.ȶ�^�Ѭ�:ÛP8�8]qy�K�l�v�$���=�M�F�'�l}��
3�~}��ҋ�C9*���Ը��c�DIͲ�q����S�lgP��_ԒhZ��=aK�� I�[���ך<�8Y��+g��K��I���'3��R2�>o�����q)��\�sb�cKJar3.�l9��S��W9�X��������ū���#�,f��ל��\��U�1f6���X�1̖�K.SSA~� ����㰆N�y޾z���[�+�#�C�&"��:�E}Ң�/Op�@=�8A^��㘓��Bj4�t3ή>�7[?cl�8E�A���'��܃�[��ޗ�9��Q�o��a���Ky����#�yhi���BO��*]0c�ځ"���/D\s��ۼ��&����(�%]dѫ����o߷7����9\Q��B���
�r��~�.���~��1��ⷍox��$�E�2�t���__8���̖1å��2<�l�d�f�S9a�s*��+x��aޗx��y�B�O�,���+�֙ԫD�v��J_�!�嚞�9���##���ʌ���x[��m��v�c�~�C_�d���s���$rd]	i�ҹd$��om;2���	�q��2�o*��K��N�t�������r`��WȯܫT������ff��o�Ӌ3�d�6�e`H���/�&w�V���Tyoj��ì����ִ�]o�78�j6�t8L���}�M��B�W�zV�5��2y��d�O0��/�oJ�8jIf��W$�Pw��h��ŀ��ac��J��įE�x��6��ʲ�9vO_+�Ɩ{N�ו�Z��/}2c �����Ȫl��;'��-�3�b�aӐ^�#�1ͥA��]�.����*.<QT���|Pi{���?*��