��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_���\Qܱ��p���	������[b-���[�������*"�q�sP�]S=ަS�[�t����}�ă��n�A��a��N1�3$4m�z|05R֔���(�鐫�a� ��?V�Lk�EZ/������%F
����ӕ�S�����ESÍ0E���u7	�#׆<���j~ \���ַX5<��"@��4�Cr�����{�R3��!�-�B�y��z���z=�,����D&"�W��g`�a�k��l����-�Dv��yR�&��VG����Or2� ���0���*;[4,��� _��}�E�C� �%K��`ڱʨXl���U��=,��oCO^�.^0C����ȋ`��,�w;ٚ�$�1ƙ۹�2us��������1���6|�-��;�6�x�o��4L�܇�:��!��g�@�����OT6�$�OZq_��=�,c��ܗ�U(V=���
B��r��<iI�i��uɅ�,���ECv��>��|�bV�Fs��_��xך�gZ��'27|��M��/I\��Yo� t�h�fp�ſ/�d����=|01r�q�[�	�K(I@�����.dt5������2n��6<�^��p+���0z2x��O�`Ր���E�ۮfOx$hw��"|b톤$!�2��8����
hݷ�͖EA��GW�Cw���:`u*���r��ڏ
��#�_@ЦΙ�g3zeϻ��v��^9p=�B/NI�5$�C�t��2�)���13��<��Pd�u����~�0ioy�˪�����3��f�,#ѭ��.�o�H�wc��r:���s��Y�����f:Q\s�ǣεVw�ɢ=�9��0�#+�tn��N��W\�����Y�����j�I�w��|_��g�����:�Y���Ŝ�����,�)�g=�i~�V�݂��ߋP���{�e �~�سI�T�N��2�6k!B�(�̞.�K{/w4�Y_x0#��1	���]�E���Q�y/�s<-vwKH4>��Q'�J�<U��S��F���Eìxt�!��u ��j����͝P�O�1�t�@���}<B8����L>\�Vg_<��ن��{��[�c�´��q�����H��ʿ0P��mc��Ce<ROf�SBBI'k��g_�xR;�	�E]�&����A�~q�����W܀oq��:�Ѹ�AT�V��b/6�Hj_0\�&�lt�?��xD��2,��G�7�?�B?&��v"�O��"&*�/��h�(�� ����sP)�eg7�-�i��&�h�m`>����ȸIK�
�4 �t�����L�Պb���_��lIBD�iphOߌ���C�H����I"�I��(�$/+rkl�~�6�c��k�^�a=E�X,Tb�t�� ?��F�^⳥K����y#�i0v�j2ș4�J#���x���k6�=1o��q�e3���n!�y'<�'T�ղ} k��
D|�����Ih"&�>���f�5w�wg����7��/��JsZ���\!�Sṥ�gN��V�@���v��>>\��-Oĩ`*P��&����P7�3�g�ێ�l�V0`�P
��s�n#��V3�*� �0�SMu��2���(��J��̄CT"�Xظ��H|+��~���7`�UR��g�a'AXd\�B��\4�	� ��$vӒ��z(���~�#P�S�6�z ��x~Q��+6x
�+��rᕶP1~�v")~	`*�3t��'�IXPUE���yKa6�c�`)�R�ա���ܧ��J~ �72	"��Ox	7�3�6��	P��bF�0�@�n+�T�	ҸE�Z{�1^$iT&+ȐJ+���4��~�o��q���n/��l�e18�|���l��c��"��&���@�d�ͥ������i �z��f�Ԕy�dN����zJc0�"�+�+}_�N�^������-�Lr�ah�+nϴ�S��d^ȝ6��ϛ��b�SL@%�j�ک{��@���J� P�0��?�B�*�o=��ϔ�9Q{��� �)�vUHFe�㰵��i�E0��x�򑰧���W�|Ӷ8,K��p���&�]�$.6�x�N#�y={Yl��tˬbJ��Cʃ�6����B��;�=�J�R��gb}�d3�! ��u�ߕ��*��eF�d+�X�?�%3	�P��͐����8|�H����ʇ���SQ5>4y�����Շ?L�\*b��q�L��j(��r�PQ*Q�����e��}k���n_I�u=5�i~M.GhbX�4V[�#QHs�J}� 7�G���"��d��dt8ț�@�C��D��J�'it��`y�T�m��~��8��8 &�k���6�j�3#��L�e"^/��$�
ͣ�f�s���r���=��zU� �������А�q>�����j��P�ɫ��2�| �~�B^Ӳa��_ٵ_�
�G24/�}f��S��4�<WӺ�@���^�o�-%V2�2W����6�➦t��x|Xh̺y䶶U�&[�@���(8��� �]NZh��s�9��-��-�r�ui\f��+=���V*t+>5��;��Q�������i�&~`y���!�WX��R��w:^����H�� ��:�����:pj�p����ĔFXf�+KQ�����c���b��˔øY�$B���B-�vx�(AThZ�}����U��\G�	���w���l˟���i8X�:�����@�s��G����,}+��"X��fX�D�<�1=e�_�&��LV�{.'mV�]R��à������iTc?�.�0�&j��x��u�bZku��&����/�e�n3����7�Ǔ�OmW۞#���qTm� c���ԃ�ם�����֙^\^Ϗ�>SC�à��d���P��n�i��ވ	�(?Jyִ!�`� %����BGp�{���y[S%��	c��0Lh<�&�jrJ"9r�����4����d嗓�ޱ���=Rz/�.�{�
(�nuV���2�h��9�	ѫ
Ľ~R3��(	����;�f�Ey�ýg���޾�=L����!Iד����7���l&��`�h�*iJ��#�1�U�OǟG��ҩ�`��អPF/_�3�u`#��_�"�%(Pyy�ʁc�ĸ��|���Ƶ��C5���2q߄�i�7q�[�ڲ#n�,ƨ�X�/yф�@
�0I�K�K�w�w��{c��lc��7���s��bۙ��/Ӥ9������6]�������Js����$f�袠�
;S�r^��"�8�G�D�a���R��/�t�u6F��%Ծg���������3I�l^�}�������Rwt/�5֋�-��?��P�A��x���!�V��w��7�.���w̜%���%�q��
y��å?����暑��I���=�<�)�":�O8h�*3a~�T��V�P���Ȕ�<S�l��hR�#��;f�i	�l�ÄB��k	rt�M�&�9��J�|F �I�n��V<*^�ӡ�u.��ү���~k('�tE�y]��,#�،ŭ�$�(����f%��Nu�R���}���]��GV"�P�mp�Ꙗ���Ai�
��ϕ(A�'~���/7�/� �M�EV��eKm혧�1z߼:|�����K|.f��E{1����][������(���cN�6VOr��I�lS%����x27��|�J�oQ���?���ym���K�2�8'�A�M�)��X%A��n?d�'5�b|�����h�Y<�q����������WG��èy�A�Y`ےU�~Z�e��@��B��{X9�s�	Rz�mj\e\ى_�F�/D��֎��`9�*c������W��3;�`ʾꑏ�vN pL!N��,X>�<o3��mƢ���>h��xI����{I(]�LB��$;�l�mt?��}nͦa5������'��-�'%ɨ��&���١�\A��] w	 �-�a�Ż�\�Z�m	ie�j��4�^*�Fބ>2�*��)�H�M�㫛�b>��}F�6�S��?�Y7�M��Uu֯��"�Z�,�L��~�UZq�����o�*̐�%��4��ɪ�����$ҁ����m���?$�ͅ�A�X�f'Cr{.D��d\:z1�w*�㤏({[�=��`-�1�m~����@��e&-��f����5��1���Z�#�M!�����]yx#l�I�+�O��s�c�v�ĥ8�X\�{ �͎�����)���C>x�?�}բ#�J�����N1��P��d}��PKbҹ�W�_�
C���Y�j	��-�O��/�g��b�&n�*'w{Ǥ*X���Lr3A�T�QIV��gc�k����*��������):o���H���¶�d
]*����p��ח�U��������7a��d�LfI��xv��4�7��|V���e<<V�*�v�!0�A������$Ŭ7U�؎���'\����-�-Z�vNM�S��kef=8�ل�ei��n�o�$�B����Gu�����B���_���]ڼ����E/�ty��T��B��m�p�s`aI"0�ѓ��o�X@�13�L����W� v�9�YY�2�
�^����F9]�L�q�v�j�Y�>��C]�K�!2ok�_ MA�D�Q|�tK��2ta��5�T/²<���	I74_�>Z�n-z����{�S)X��^ ��W'��p�����`ɠ۰�����|�(��HƩD�Ա�/����Z��%���W
5	E�u�H�Z����ws	��˖��r�mEWO3"��w�3���ہ�����v����X�!}k�s��'i�M�H?ҭ�d�r;s|sR�jr�u���v|�ނJ:�J�oy] ��}��<m�4������g��ϔ�`[��T~�w�?����Vg�Q׻3�K#<N�c���{0������s�3w�}��{~�u(c��l$��%FXj`(��dWy�=tV��.����kӓ{�q�C���n�'�hD�p�Ԧ9an�K}�O~��荢� u�t�:��m��,��6�?&�n �pq�㬺W��e����]f����Zl��-��Dr�DO��'
b�/��E�?�Κ*̡x���kuYN�֪�r�!;$�9�(/�m��r��O������L���b�͟�ǫ�n���o�႔���5%�{�����Ѷ�{$�b����)�ئ,�o'��t�n	��:Ef��Ny&s�I���eA���ݳ�e�:k4���q�n�,�TS�Iݥ})��˓�Q��{��\\7��+w����:=	$1��şԩ;�7�z轲X���3��	��4�}� ��W��g�0�ˋ����o4ݰ6�V��c�_����پ~�89�⛎��D(Em�<_���&%v����=3����?<q	�,0�P�E��U	73�J��x�t8 lj�Uq7[c��oZ.'1�����A/��Xi��V��W�gy1�����i�_Lͳa���D���~=�4��V��F@�����V�~�轻�L��#�J\Z����i2�}vK"�]s��5ՙq���|� WGj���}W#j���&a`�'��M�-,[��7�f��u^�E�����Z��R=&
��{�,Gi�i��O&�Yz>q��<��EIyQt��a
��2h;�_��"��l����y�����j�-��"	�B�Su*�F%�eZ��\�~ti�l(��˞3�g�f	���o�k3�L���qH�N�͐` �P���R@���`��.����ث̤���W����b[;���q�^����b����,�6x�s�/�@3�R�g\BɁ��]�,^|)������r�P"�=X�O�|���=��6װѫ�$(t>�6��e�R�|tt�7��"�#篘zT�r/Z)~A\,�~����:����*;QM5����gy�3w,4r��wBh��OJJ�0����eC7֥���HVd��G-��5γ�f��dȪo�B�T:��ʱ\~cR�0N�;��M�E��%�]��[-�q����lKRS������Y�8:s]�3��,���=5a�9l.���[ ��,ou䶶]�H�#���i���$61ԉ��b�R���`��{���4�^|G)PYx&`@qw`� �e���o쬛����ӑ��������rT���x��M�z&zn��`��^3���	�/P����#}L˯;��@q�a�U��&�=Z�uD�ô*$�������Ex��#Ǘi����F�Ȳ)~�w�1���oF�����,N�j�O��k3��,}S_7�ikzs��Nk�R$�LY�E��w����|p�Fg%��RL)�K����&��E��V���"J�U�ѷw�@�v\��dWqI��ǳ~��:;&VR�b�h4��G���o���Mй���]� ȝ�����1�6;"Hlf6�\.Ģ�
���ewS��u����t�Vx��2b36*�g����.U%�m*.�H���3�h/�����ڗ�S
\�����E]m J�X֮�u��]l:�x]u��V5��IX�W�rߩ�|���}�)#!����y�G�� lZt;y���`�cj����C�젖�9�b{t�3�Q\�xc�'�6
Uk(G�%�C䟴�?_�m���km����rp�/��,�X�&�7zAX=�lQD��䇳ݽ.ԁ���t'�ª�s�J5��-T����vyh�c����O����5;���b-h���o���RP9�{����؉=��Y@����ؓ��6SK�$�ڒ{;�kC���GoY��a�D��=_�t:l���q�'���y7����+��Y���b� ?y�z���	ŵ�G|&�Q�)�*u���/���������~�f+Q��־�Iy]�j��BbO4�!j�m��3�.߁j���h#�����9%�(��w�׫����ϵ��6����%���m�`�iUS�?k����.��}�e��q���J�������B5*M��F��c��ؒR5#n����#���nM�ԙ��(�9X���ަF�.�Fnz�H����1j=��R���+nc7&��kVC㕍�ٖ��L����gɥ�"fZHV<��V�����e{oĜ���H��A���ґx���;zAk�a����J�T�Z���-ݧ7���{��N�>n�3��ּ�(Ҥp&]�Ø�տ�K�o9����zn:��W:�O�j����1\��N�U�,�<�t�SB朼Z>�b��.�#D����
�<V*Ȝ���sM�i�F�\��n6[?	]��/����WS!.�(�!<D��?���ę_ھGN`���k��:�X��	$���ڿ��^%�5��(p!��"�:����~l�$��Zۤ62�W��j;7+�q]r�W���u�͋��'>��|��9�YQ���ʴO���^'�0��<��i~Fjӊ��H���6]�&�؝t<�F?�l�?B,�|��>"�O �1E���Ȑ��U&�,�V����^�-v���\��@�1y���G5���QI�o�.�)xrHH�_'A�����B��ǭC��C)��9��`���Y7"<4v��f�q�NYC_�|�Ǿ��(�9#h`́�#jB�Q���sz
+u4��7
����
Fd�$�o��%f�R��!�nH��e�9�Z���g=+��^٦)��@�2p`e׀�] S�|"���JF�=M�:e5�')��}��,�͟��Ji��/jy�9����K8�s���L��5�@K4�{�Xh�e�����l^�Nx�%~t\�JH��n�Cu*�9+�����+(r��M�=���e���$�b�I�1Pjy�|����[Jq+��ݝq��i.���K�'t�~D�)C�bsǒ�4��G�zPٿ�~ES�)��,�'��|$3G�����
�Sm�w;@Zx�h��/��$ W�y?�N���'u��>���>V�c��C�jݛTz���A����g�:�\��v����O��EZؘ��CQQ(.h��Ђ�S�3w��-}���Z
���<��.3hc(U$g�3x@��i��5��ڱ����+�{ZH�|6�H4uv%�V8A���,�r���L�A�&#�13��j������?�!�}�9rce2c_Ü�9���+�`n�aB���i� �,����iA���mxm�_R�؊!�KȿpI#ca��0�6$S;�UM)H)���ͧ���j'�ᔷ����A�*�H 0ER[����rU�?��Y��U Qk����R�&��!���
}�*�1��"��wj�>��E���G^׌��|��qW��~�y�>V��;p���U�D`W٦��3��@͉;N@,��ۏ⡏�R
C�1N?TF?r�Ǉ���%��"Q�K�w��ceoh�&�`�i��������Q��J�f��E�L4�w/:��	��G�'7�ѧ�������TXX�I��iw*���D:����I�D��m��قM�m7�/�y��I����5�Q����/dY��PeҐ���׎����]�:z&�H9�����Y���S��K�ӷ�8 E�~1:�2*���(�C���F�#t9@�;���+P�wB�m���1�m�a���A�J�<-�I��#.�Z7�
y��ʀ�t5����>��R���U����7�����m(��YcV�ӱ�fJ�|���kn�)b�}0
�|m�ϻ�/RHt��Z<�A$�z����Z0�
��䪡�eoCv�\�|~�0�St��a��p暠�h�ǍrsyA1���e�x&"D.�ݴ����f�P����P� �4N�q�u�ϲ�^�R��4�o� ѴÔG�(K�'�a�sp��ޕD (�)�i��DV�H �z-%�F�L-Xұ�Ց�gtRI�Ptk�S m�r�bj��|؅�`����5H6�J��;�;�XB�w|������iRG 5�m(V��2���M�R�χ�=�R��\�b*�d�4X�4Z���"S��Tw�3��yi�׽�����x���A�q]�[�|����cF�\��;E�
Ac�0�[֕D[ӥjBG�����SE�v,(5D�-�{�ڠ�sj�
�{��� 9/�T��&�t�8��[��&~����Ep�19�䓥�5 E*�Zȕ��_}ͽ�=��uZMc��v��#�X��b/�������pFR4�=j����1j�ORUښ��KaЎ;S
�'��XN�dʖث"�|/G�Rn�ڋ�?��2��COj�qz̥qho��wn�Lwo�'�ֱ��A�E1Z�E,n�����DE�7��tP��
�}�Q1���r;���9��g����:ݰ9�d���ӓ��&�'Am�<}MBʾ|ć�df!� :���/P臙�8$e�X[���Ů�VBN��J������n3̳�D�3Y��}�R�Ul�+��W<��<R2�e�k�CK�Ņ�|~���pj��#z��#�_`�(w�UKs��VG�(��
�<��x#�:���8U�n�9�#W���2v�zY��M�i��ٻ�Q�t�H�s))0���$K�Y���K�%*I��Z�2S^nN�]���*�04��F8��ǫrGn!${Ә6}�P��+�g'y!��Յk��tG.]Pvw�������[Պ�@I.�G���0�<���`>�\���Nk�¦ʸ�|36Pu炰a"kUap�6��1�#�,O��nQ����t~�i�����KE��^x���?�*m��/����f�/�������"�^nus����RKq[ �c�V���6�`\m,�!jz�G+�q�W"W�F��ų��%|Hb�F:�Q�O$�g�$�*E�`��n�M�m% ���DY+S_o�Y%����aM�`�&:�N����N�X�8���������j�#��1��H؇"�����z���J������ѵśQ7!�̓�u(E�O|4�쪃�4+���l�.�Js޴�����v~�9�b("��� ĵ�꽇��(]A�	M�~� �9���\[u}�]E��݃��s�%+�Ϟ2�X�lݎA��}�ꍏ�1l\�.ۣXބw��>�,&,w�p�>�����o����)S�>��''x��V��9D�{�׺�J��������|�-�z��8Z����D��]�L�,�G}W�d����}���xI`ܫ�z
=(��c�׍�h����b�"�{��c�!Ϧw�q�E��8o��ͮ�<�tx7:mn���.�/0)��e���e	�l�2�����^teR��1�K�U�I"�_3e�~¿����mm��$h~��|�/�$�gn��vl��]��I�w��v&U(��Z�ю�h���q�B/��������aBz�FV���삶�a$�>�ּ�Q^��j�/?\����m�^/���qP�I���&񄤋%;��%61�7��WO�EAeҲ�b�i��X��aIob�
`w�u�+��gw�>zق�����e�c�@H�H��1�T�J� �ͣMřMqA�|˭UDIj'�H�L�H����N���UO.h�?����P^FUס$`�~��Ц1-�nQ�a7d�}�:�-�g��Mv'?�i�j����g����E�O�N�#Ɍ�1i�a1Lh��_���ꯌ�y@dG`	��Z��K#d����?��uPTX^GK*�4�n�w2���ǖ<ؘQ�g���'=U�Ȝ�bȵ���"$i* ��*�އw�	j��2~>��]���t�����c�H��S"�%�Պ��9Yƫ�շ�����3ί;$`�K=g�r��P��+�����!��ŷ���Y��t��'��d��j��P��>Z�B�d��;f�l��N.�^�>�p�qWm!8�3���x|>1?(dF����Q`re/eUT鞖n��<��q;��nf�q��Gb(�|mO���G� yl��|5��2����	ެ�⼴yQ2�����<�Y�_�W�ga���F��<�O��D1��/4��Ҩp��_[�p��^D�I��R�}���(�f5�Ѧ�+�s�n��
�jj!�����|�ϰ(�ͩH>�M��i]�N��Ӳ�7��$9��k�~z��;���S�/K~��Jr�K���
�L� ��L#�'�b��X��C���I���h��KX���-j�6�����;�(>��@��n��%�&��z�qõb�l��C� }l��ˬ�[l����̕�}|Tc-������@	�Rp�Ƣ|�l���+ݧ��>��H#向<���t�V��k�h��z����Fr/��!�+��h�!�Q+[L��Kz�,����~����uY��V�4�0�;Z�jE�dy���5oy���4%^)o-��5����;Z��0�U<��{��p��Z^�[�T�L#|��M�~�m}i��XRE+�3i����������D,鎶O�*����Oǋ�8�����˩�}a�j��+�*��b2����$��n�cv+��5%`�E7Y]=c�g�3��b�y��K�e��+�`Р~�˗g��z�ڎE�\&5��Of����	�Lƍ������TL��e� �h��ۑ����%t�^s|������z2���p�٘��f@�$�"g�A��zv6Ƥ�E�T���PJ�A����l���6���Q������:�-�2P��
eif�M�n���(7�e��g%ƣ�+�8�£#-D��2y�vRu���/����	j��3��AaA{��[����X����rij��X��-�q���?(,W�գY�Vж"a��~L�fA	�8 >~��V�_�m�����DM.�ߒ�?��v3U�ٽ�Vm��F� �c�D
����!�Q�I�٬1!�I����`���,/A���v�E��Oi��t*�!�����J0�μ�r���eo�ȩ��zhL�U���:$Z��s�ѵ��\�JC�䢪�P�E��GL������-;n���\d���2,R/RC��D�I��*�H���7�pN�%UZ"�+cX<>����5���"?�id��2�Fڹn��c+��A��[�Y�D�F��a��f�%n��asr�XvQ�i-}VU�ܪ���L6ٚ5,-��W4l9ͯ���,�����2XX�e8S*�h`Ep�t���?�!j�ru�Ex�?y��V$�[�3C�����a�pD�VLn�v��?���b�b�v��fni(rݬO$��.h�^"���B+�����#)ꦀ>Ƥ1�bf�֥Ԗ ��螚��Rڞ #F���YK��r�14���&��2�e���{�x�Ձ&�\�9UNV^(��_.f���Y����+b�Ñ��f��G\��_�-���Y��iG�_�C�7�����5	��L��qCw�U�MS%�i�:{��vQ�/���N�)�mk�������rR�I�
�O��
&����&،���3��mE>
���X�O��>]*�ЦN����v8���o�5χ׺(�d�=���T��*�rfh�o� sN(}��1��G�z�M� ���GI�x�����K��A�����.���$"4b����̜i��x��4�,	���չ���_��*Q�L(?�{M��u��"����[&U�C�9�Pb|6N��t@Bo���%�N�3���VH��5�(�Eku�+H,Z�1�� �u8��P'ztt�$�;�w��4��Q�����]l�̩�:+Ȅ���e��a����L@P�7CB��ME�DL����|g�K���"�*a�B�^���O�AcP,)�ao��n���c��Ltە��j��U�}�+m-�靕�5@:Z���c�~h�$DB17�~Ǝ7��J�}`��5��hmQ۝�
�^��Q��o�T��-��>y��I�e
x�;����S����P��{]�!'_����ռ�n5������D�%�i����S&�����bS��WC꒞��beA]h�r4g){��^�E�3�u[�J�v��Z��9�H`<�lĴ��ph�=���>}�)�(��������3�)zl�N�cwf��f�5�����0�mQl��,s+̧�$h^7"�!��]��|&����v��C��8�3 ⾣�
��/�����M%�"����{ �ܡ��q�� �)W}Dn��.Q�������CF�1�d�,�>U���D��]�k޳;:�2����L��d�e��8����RE*j�7�݊��.ʝ��"G�q�6����;���G���5�l�P1��c�]4���+q
-j�3w(������d���)��d�ْT�V�t�X��P������T�ϡx�s������#$-{�z���ď��~���x��	�/zQ�t��m7�^wE>)���R���&e����Ǜ;^�x���9`��>�{�	�O�58�,���- ����N���	z�%�G�2h�}b��s7�,�Ϻ���k�/]l��^e��r�4@u����~s��{�9,�VU��Wð����.P���B�I��]h���e�t<��դ�0�͓�h�[ܮ��G��Z��[�:h�H?�g��@�®���q0<��k�%�U�������h�I*�oZ�TB:k�$��y+ 2�&��7%�U���?1Mw���0RیӃܵ�*l�l
W�VZ���r���#�Tϫ���n�'��!��{�BW-N��D�K0WvR�H�O�q�����}Cy�[��)!x�=Pvd�&��"+��{���?�M.��#������nzR���0F���ņ^�6i��%~�R
��-�S����v����u��o`=ɅG��g~i��ڔ�'F�j��+���%�2�u�}�ڭ4��k;Sj{��%W�Q��o�Bm��>yp��p�����i�DZ�� [W?�Ԯ)�� ��i4�G�Bw�(=u�����G�e�zW��cH��X�+4�$1���7saX)���D�����~u[U�{�N��]�Y1��D��E��wֲ�~�9�7-w�!B�S#2�i������*��/,Yl��N��'i��c����U��)	�q��'
fN��~����z������+�T���c	�V.�돥���G9|;a(���A�v:�Rl�'���]g�F� T4y_\v��kxM�@����,�V�NW�	���@$q�y]����t)?��G�$0u�54K��Y����Y�[�l����{��`K>x�fz�	����e���}��8 +َ͘�w�z��n��=��	�t �7$0��%�n�n ����`��Q�\MX�eUٹ�|���T4��ǐ#���PG僊���h���-�r�Z�l�9P��+6A����1"8Z:j� 7��d���<�o���tcG��j��ӱڶx��ӣ.,��,\�/����l߹��:$|=?�G�E�;nQ��u���'�[�؀�������|�^qP�y������%3懂�-㛰�6�Hʹ��`�~?��sv/��V�E�7�2����=S�z`���Qr�� �#�ģY���ڽ�Z�;G�v-i���ٖ���*�̈AIaH�o�fW��;!�r�sRX,��$u�k��QH�og���z&~��GzW6�-v�p��=,[ h���7P�CQcx�|�����~R�?\���hBv�	ܐ6��[��2r�k�Ui��<N�n����w�����s��y�h�GV�l.:����E��q��'��!�\��p�~�� �Z���`?�`����T�;T[�K�=?�*
����-��+�E�ɇ�S�qV��?�=��e�
⢍9S�16P��W��u��\׺<%VD�ŉx��{~���`FT�8�^P0��ڬ8[�����p;����,;��D1��-'m;c���G������+�+<�X����_6]�|ө��+yY^��U,{�������ǡ
w���=R`��Ӹ�p{��<��ޔ��7�_�W,�F���j=XֽMP���v���� `��z���v^2�ߩ��hW߱�����V��C��ӿ�T��3$B��i� o�Z8���~���_�TAR�"s`�aB+���.5�@���&@4���Z�Jַ���C�'��"I���	1��7��BS2xt��,,��.�v��m��q�!��"?4�'v�W��E?�-��];܏1�b�EJ�b�����qC�e�����P���|�(Ѱ����!��"�z�AU���otm[4��."�`�W��f�#o-�G7L��R�/�h�O�RL��q�v����8YY�%�3�(�4n�(A�J�Λ������
��}-7����og��3�$X����^�_�Q��E��vs�U�v��hʞ6Ů��h�?qz�JA��a�c�����	1?>�O����^�c�c?��1�'Q ے��R�Fa�:n5B|]��Q2��[�@r7���A�9����F�ӓL��:F�^�����Է�S0w�Ӕ���<ϕk��s��K��4�#�����O�����H$�B,p�]9+X(pp���-���<�aP!fw�Y�x���`�327�2��3oz�׳K�6�tr�'�w��Ӟ��$Ci��g��.���Q���F���V�BSa��Q��u8��7���p�`���lZ����� �����iU^����P@�Q:�K���J��H����ń�^⍘b�f�u���/^����+�|Ի n��Q&�g�]��TXgu��j��d��&q�(s�p�~2�_<	$�mL�X����VK����g��@�:���b(�P�Zsjx���b.�E��2����	:	����C���lO�OY�CUj��#ًU��cR�X
P�۲�"�b{y��T^.�2�p��p�(L��++����V"y���qJF���!a���I�Db�=��[(a��!`�P�/���$ys�n;�%(� Z|y(�U����/���TZ3ɮ� �i��M2���'
�r��:5���v|�.���+|�;�d���>��N�iP1�f�Y��8g�~���K��Nԯ�ōޗj����3����Vj�'�Z\��Nl>���!Ӄ���6 ��i+kޕ����>�E�d]��!���S�V��́��{� ��9��θr�ɦ݇mD��H�6���N�^!㻳c��]ɓ���H���8H����>�9�&����S����ݳ}PA>7�L0��8�Aԁ#��;4$���Y��v�9V颓�_-�9�T�6	vU)ĠÝ;-����fiL�3G��6�g�[�Z��� �<$q.	{��"N0��%+��/dO?�¤f����F�@�JP�����;��3q��a]��3��Yp�|_%Ў�ݫ+�NY�GC�t+�}-��ٛ���F�ϣ=a�6w��ߩ?������� �W�42�r8�>�MM����&4�a+v��+{+Q-�5�4X/�k�֑2�l���NR���i�"�-�pJ9�p�Y��ā���w�+r��f��'&����0��p2T+(�j�6��E%D\��k��om�["�l��F�������O�t��ֲ��p-��ndD�������.gA���Y�j2We/���g�zuF�zw��OᭁㆯQ��z�-�����'�p��g�Q�o�f��*��Ԃ��_�jG����M���"�	w���s�i}CL<0���=��]*F(�./I}�r �S5���HSQ�x�<-�xz��&�1t�������V��6��E��jPΌ��]�Ǟ����V�zv�!'���x��A��&,�J�Au���N��l����48h�󤢍���<w_	YJ_��[C���z�W@)�D�6�pԈ�-�}Ȫ�[�/U ԩ8�S}�Tߤ��tu�s4a��l�Rtv��ֻe���<���� �
N9�Ϗ��p9��d��@�lgLպ�^��Iw>*"K �o�i�h� /���))ϛ����+ڴ��� {K�w9�"��r�� 3���t���%���μ|j��Y�='�V��������1>aM���R<�D�r ,^
4F�N`�n�!��O��7�A�����L	�g�z�iø��i���8c��@<��X�)@ҝu͠dfٮ�S�:���-ĻCB�'?8��[C��p�GXU4)5����-,���K8�����UO��g�����������\�~'���G=a�R�3s;��'�/2񵗡�K�����	��3�{� { ����Sm����@eB�$�,�E�����߆�Xh}�D}ⷨfN�Y*����p����A�H�/:����g�D]�fë�	��;mj�S��#����>M~�P�60Q�g�@�&�&5ku���3=�7H�8ܠ�S�T:H�9��v˵��$h��lx?Yjm�t�{z�R9+u|�+$ ��F�~�
]�w���?���o���U䨃{�f�i5��M��jpK[n���輱p��Bd�Qj�)3�c�H�~E�П2'�y�t��*bb��iG����,3�5����o���y�;�-�-�l�RL�^�oe;����͖��(�Kh߿_9�G�Nh�	T�O�/#�t�R�Ǐҭ^��5_%�A��HW/5f!��b���b	��Ŭu�	S½��yv�������y������9�=�[�eʂ���͞	���C�$�cѦ-Ɯ�zb�D	
���l�!a���c-ۨ��#�?���{Uq���Qk]�9�3%f��̅.V��ff?׊Jܧ��gҼ�<G �;�����7{�S��ß@4�-���U��`UN�[���3'njS���ĩ���8�� �@���|Gc4sOp5{/�ށ�*������$=Ψ�{�������bIC�F����� g������Xi0lN���f.��;F
;����
�mۭE��C��@�6�,fی�,���������ݗ����AF�kHKz��%@ܘ�Bnb��9�o,D��cp�l��ec���'�R����AH<��@TU�ԱH�|+��/VHi%V�m�=��J�Ds�|�~�OU@;�o)�AϏ�,��m�Q8vJKn�e��~(�K������#pT�%"(�#���u�;Zv�tKt����s��y`����8n�����zR��I�v�WC�� `��ZV�Nmx�Q�����	��;���#�T��h�v��?i|���'��K�{.��������"����)��p��_���m����q���J�a�by��Cd$6Ah5!H���G�E���"A-��atF!�����g�[��7�4����'\)�ʑ,������N.<��T7����9�.��ar}w��pF[��������0��x.sE�:�O�%�$o�f�i�El�*1$>�y���>��I�#c�i�Y��y|b�ue(d����$P�S^��D)�B��VwV; �\<�=f�e�T�YQ^����|&,��绞لpb���Puc��M��=�%�s~�a��4^�����<��!�Ե�tX��x�F��a����BD���vl?seЉOe��N��q�A��������ci�ǟ�	��%�[��(FN?Ҙ(k�:���%�`�Ul��y�z�a%�7�?�_sP�w����CG�k��7h�2dӻ4	�����-��nc��2ǃ�j�GeJ����0���
�j��f�>f�ז8���?���P0;Ir�6I��n��L�U�j ���z�'�7����K62���5J؎��JU<��t�Fm�Ȏ��2����wy{��@z�ᗌ?��y�ԋ8�cv�̦��ly6����M�y�#�P��i�x1f�`�دȎz���Q�E>1���'�*;�C0#L���qD�'[��cL�D+q$rO2�N���_c�!$n�0f�����f"���@VЋ&� �Z�A��^{�
ݥ�Gв2�D��l��ܭƘ���T����3=��������}Q��<(b�.d9
o9�-5Y��ކ����R�皰+ҡ�׽�f��MHB���QM�{�仲�3b��m낺z=��E{�O�1�-î"���
���  �k%����	R� 5;�E�)J5̉h�W%%S��@*��e$�5���`f�q]���?ne�oP1[�?���-��Z�g��3j%c�r��`ˎR��صh���Y�'�cS�:����f����bp�ۡ@�u%d #�W�k��o�(����43��A'��O��p��}qQKy����Nf/x �H� A���U�B�S�Ҝ��w8ԭ�|�s�2�o��2��́"%��~IZ�L����VA�f<�JAL�t��DD��'�FE�Þ0�8��T��`�}���:!q5ײ�j�ř�N�L��P��W�c`���a�-���I(!��S���r2,b���q�1�H)i�J�e-���h�:C�7b��f9�X����_	���.|�n��#�rO�_����,1�f�.���sܸI�ֲ��{e�-��^���Y�p�/�r
-X	G�����ͤ��܆�(��۪V�K��c����?��W�V�F��hP��V�2z�+��b��N?��]H��DV�`t��9#�8�H���fP~m�L��pC~*ǿZ��c�G5 ��#eN��[��EM����TX[p����0�|-�<�FJ��H�>��Q(�� �N_/W˳ك���&��-9��Qdv([��C���}&+�}��n�I��^�VZ쫔k%V�NL��a%ji�fepy�ȀE�B�i��Y#�/�3��Ÿ���yH�w_�S�\q�ɜ1	����$�w8�;>!�;�r�6>}�_LЭ�O@�[�v�z�2��1!o6�H�)ZW[|OiH7l�XI��A�H��/�${w�ݿ$̝NI	����}�b��R���T�M6ȡL�������A��u9ze=6��V\f��^\�t��-Q��������5	Nt{Gj1��->H�3	w߫�4�.$b�J��M�y���!	�S�Qg;}�|�w+�pVL�r����_�>f��`܊��(-�'���ƍ��ұ2�QM�;Ҏ���F��hL��~EH	(s��ޕ�x16���a��?�/ g�� j����?*�����1���wo���1řԧԿt��Ŧ�aC?��3�짘���+=�/��
y�t-ќ�D]-Az��Ls݆D�dx�� �5��5q,&����h�{���=;A��6��zN.��x���g㨠��4�$q*9/�b1Qc�n������u��v�>��Lq�ս�рtZ`m��>��ڛZ=��Qq��76 _��e�:(�23F����%�p/x��Ӌ�:(�	z�M�|H�dS7Z,�^g��q%G�8�iS�\�=����� �ߍެ�Pwێߢlp�M���FmR���2�i%5����OO�|s&��Q�O���f]����J��2��b�H$f���#��K�1�qW��G�N,y)vpeM���_#(9�\lV��@^%����6u��.wBf�ŵ�/Ch@�w"�?���#�װ}�Q(6�hź�٬W�ͯd'���_��?¢F{�-��p��vp;�,�5,���Ƿx �Tl�����\ز�|.�0g�/:{UJ�9����o�t������L�Ȼz���D�dha�ӑY��L�5߭`���U��b����<��\�Ö����E�z�og/{��5ŀ���X6�SLF�~��A�T�q��1��z�0�P�<�}���Xw�~ITn��X)�&S%[|����6P�Y,���k��*C�|ĒT�����$0���C>��@��N���j x�[	}�Y�qY4�� 0�-�Է�����f�:��8�ډ8+NOf$𼟵r�	�c�{r.�6(0	��~�Ȏ�ǌ�4���!B�X�Ak�X��!��BJL�D�PK��4�^Zw,��yz+׽/����<ş!l)|)I��lc��Nue*��1�n��l�@Y����d۰+������z%�-R�HbY�[P���ms��x��ԍ�d������n��]�1�P�;X������DP��k�0��)����m���Ү@9:G��5��h;$���d�! v*%T��`�A�l�q&���N�$�O������X���9;�=c.X;���Ɓ��,��=2/o����Ξ/��!�9	A���K_�±�����t#��%zgE�W��*s�QQ�Oϻ����G1c�
�ڈ׆�:2�z�0�0Cv��W��@=D���i<��ā劾֩��2�Ak7�e�';�lƶ6U9���T�4(JH��˚�8#]��qs4}���R��-)2�z勶7��Sy=���S3X�4�����{��z�Tm��'��B\ƻ#�2E�:v\�\���L����t�:�?�Sf��eZ���M0td�!�R^�e�jMR}�8�Y��7LL�ݰ���q~�O��z~N�af��i��e�H���*b�D�m������9?����]>���:�ẖ��2�W�UBT�ө:��k�-�ڼ���2W�E��_3�TC��N��gcue�i�w����(���e%����y��吳W5�/�a3^a��onbP���wU�cz՝�*�Ns��r��3�D�� A:���ϻYx��<@Y]M��Ӻ:%6�^K�X�/��4(R s�/`>��-�3	`�8�_N+Cn2s�zdH��}&<M�ߦ���a;@˨����<�Z���q�{�R�-tA�B�9�Wm	�$_��[&;QQX�#��\k�#X-���K���?�Ks"�]*<&+��"��L�B"l��,���1����Q��]��Qp|Y���*��Ҽ��'3��-=�m ����NJ����ݑ˨���+�F�o�!� 2�78�)p�������*�$�O>��o���N`1Mi1��m��<���.(j��R7�C�0�q|*G�dK�����fgL�[��</���\C+�9��{@3Ե�<Gf�N�NX�J�sE�3�������m������.K�应�뭎�-�R�UN�I�������;���:}?�HE������OYIv��.__	ȵЮ���^��@��G�TE`��-I��\��C��Z�_;TO�_#��&-�c.��O#�l�*�&G��#5�/��KZP,ހ	X�^SS������q6�����!��2?d5뱧YYǞ�P�s��X�j�c�"�hg�<�~�N[rqZ��wѸ�l6ۭ<��	Jߝ�Jmz(�v��}7ʟ�B6��A��z~���(����`��!�j��8�ٓ:f�7�/�_+ϸ���m�љȺ���&�<ϗ��
CĚ^ �������V�5��2{+{�{;rV-
�u�1�x 'c,=��91��)QH'��0�D�j�"-�pM�)�%���<�+M&G�!qt-��`wʩ�_�7��2�d�;A��8pviQ��oJ2 .B����w�`�wX�����YX D�E�J�y�G*���)l(�У�-�2v�'P�(q�9te+� ]�UcW �q��Ǣ���y�Ǯߙ��\a)�OD�V�9�"�l^���Æ�9�h��9E����)οe��$�~:�L�W�n�c{c�a���f<��`�4�H�ī�9з��#��2�\��`l�)�l�L~��Fyɸ5 ��R�o֊u�ń�U���4Ϝ|02[Pn�^}�S`8��{?�0tF:&ESn�ݳeվ�)ym�)4�h�D�D�XG��K��l�=&����SvOCrIu[����zc\���؁}�S�IA��彛)�K{ixi�%9$h��/���I�l(];;@@�[��*]�E(�~���l�
�'&�-.�����Q^_OLRQ����v���/O)AE���Icyvv%��u��E3��6���Hm=^{��c��X��uُ.a�����$�iEBmy�3b���*����7K�r���"���+��}�H�����\��1^�_7ǸڽLŻ������v��@#Ȟ�X@/=�g[_��<ߛ�X��̞,��/Z%��f�x��s�w��D��8s��p��4̵l:��rХs
��ǃ�b"�H�(D����\��֌ė��:<��0�gr8^*T�!ɳΎ���\;�лjh9F�e�
��*�����x�aL�F��7V�; �{�̾�;��U(�菄}��w�gKC�&�����GȚ�A��x����k��7�<mg�Ls���#���-P!G.�l��p��暾V���'�ry�p��� �)�_ܖHJ����\Bșw/�ON�N�� זN��n��P�RCB��O_)(ޘ�َ[@୳whݷ�;\u<��f���s�fث�H�$��[U��g ��JdP ,��C�@����g~m+K΂-����V`�
R����j�˰t2����e�<� �--��vT�	�6c@Ĵ���/O���Bc�3���z�	�D]H����Ҥ�r�<��9,�a|a���lm[O6�b=�d�r�y7:EH�+�6g�)���DM�9>�I�#,���ȇ\@�u;[���K��T��-����~�gޫk ܈ÿu�A1U��H�Ӳb�W"(O�"ꂲ�r�����pqƊ��D�m�bg�jZ�cӚ����>�?���Ԗ��(��wr�C�u��Y������oo8p.(������ w�$rjkw��y��n�5��;`e�b�i��8�`��6�g}���mzD�q�gX$��H)��#��vZQ�����YPȯ0����#�#�{v.�ă�ي��cWR�j�ux嘈�4+�Y��-��n���z�8voW�K�6�L��圇V/�H	%ţ�������Lp2<NȻ�E��u쉰=I!�y9��c���m�j>� ������ {pݹy���W��<�o��4U�z�f�ynX�s"�<)���5���6j@���wyz�d�l��r�5L�)����>��ƕ��ˈ��힆��0���U(%,?{3Hz��һE'��%E�'���~M��Aʰ����b6�7�%�/bq�6ƚUl̔�Љ�E�O�`_�9]Q�r�Y�������|E\�����.��|�3?�������3hO$�nd�[�}vQ��G����>C�K����?���(b#�4;PL���}���}��r,�����x��(f��y�c�� �m;�j�2#-�Nz�A-���̲T@��Y�����#�U�Bs��*C9I�(g#e^Mdw�Tq�{��}�,%t�؆��<�6�ߌ/_ZS7�9���{���}~}���U��-�Qtjf/��x�Z�	�U<Aֈc,��Ci`��s��7�zY�B�T�<�>�7*ݚ	ȡ6�p�#������I;�mP��;l���hMے��P���v�僉��Qn��Kd@HoS�.<��X�U���p���;�׌enE�l ��,�56!��k�v����>�!�x�- �ڭ������L�G���O]��Ѕ�O�3f���������,Y<�|��I��t$��񁰀j)��i8b�`p)2�zEI��Cd�JW�bV�n�$7���od�P��v@d�H�8<q��E���j�HZ|uJ�g��K�Y��8�j�5��ہ���X��L�emn��]�X�uYt�TD�zI�H�i��-/��z��4��6��1�jD�?P��8��}�э�ݥ"f\2�q����pI�)�T�O���z�����?�I[����%B�=d���i���n�#/�3G˂���Wc]�u��ȷ��@�`@�j�窓H�)9�9�����B4;�BH�~g��ƀ
+�v��cu�Km�Ld��Y{��l#ratr�'����qQA|��۽x̛�_ڞ!{���e��Unp»;
y�ǭ[�h�[[1�v��v;GƟ"�Y[/}���il<�����9�DA��q�i��Q�M����_��h������
��%z�3�@�+9<D]��|���Ssc͜�n�6f�"���Lz�	7fh���s̛��F*i�!X��/tVOZD.������ػw`V��c-��{4�AXyc�>̅iSv.s���JUns���g>�n$?\R��٘�`����{���+���=�1@���\���hC�m��T0/�s��ػ�w
)&�g���M(-�(|O��H�Q,�ka9�����f�a!y\Gqz�i9�Ă��D�V��:��!?� �4�rC�9f�d�^����$1��s�r�4x�)��.ҭ���eK�|�U�|)� Z)��I}��;��{x�����A� �R�u�e�9�ϥ>��w��[�Ҕ��`��q�-A�r	�M!����7QN�?�y,��bm�2�^�j��ɠ��a?�{O^���+��L%-�g��	4���<~�:�g���j�L�J�N))����H����-{�#�K�cS�]O��m� G�=�~���Cl��s�l �N(e]$����*l�D2���6�f����#��6�v�!o���؇���VU`�כN����\���Յ
�U��D�Y'hz1X��NFg{v���,ZD_�?��$I;f�]dN�#��{���X?*g.+5�p®S^���w�3����'��ߠ��|�tЭ|������@7���]�$r�Lk�L�\�?�,Ǉ����b]��G��ݘ���P�fX������U�~��3(�p�)ڑ`b��&6�F2=1�u����/U�H�.�S�HM��F�U���p(N�Q ����b���֣���h���[B��k���d�+�&A�STo̮��t$�y��Ӡ}�`�tz��لJ�<-�����vQ̛�a���wJKy���G�� ��*D�E����
a�k���MBV� ���ۧgx��]]|��/�YId���j[��2!Yi+�"��[C�-{0$�a����D�ŏ��c��Htz<��K����RB���� 6�)ƠW���x�Kj��w�0�b.��B��qՔ��e�(�}��z=]����	�?2S���{|T�!�:"k9r���K6Q0w�d��W%,��Q�46ΔaW"� �������;���S�B?��J?Q�X�~�,�ï�^%�#ţ�/0~	FX��u�N�݈i�_b-�?/����/�<���q_~�*wfvu81ڳ�`k��������\lMF���HrpӴ�W\jU%|T��\Z~Z��aj���}��EfR�w��g2�"`��>�m�5�m�ω������Q�ۓ��9�����^�� Z��m�D���,���a�	[[4����o�mX���U��q�(n�HSN4�0� �kQ[R�pڎ��,��\�J��k\|�vہ���* E�]F⭛!�� 5�dz&��˶�E嵎)!�7qȄ��m��WxW���L��`����|K)��+���>�c���i�Un�E�DP�7
[z�����w;E�����r5E�D��+	�y98B@���7	���MFKM_�U�9+�R�=&O�/����c��'�y��T�vkH���t.��e�^��I9}��6��!��s;0��n̆�6�'���]?����!���ȱo:�ű�r��.ʇ��y�w�tt٠���l)��X"^�=�d����q�G"S��t|�B��}��A��M��RG�"�c�bv��k�)
�{�wu%�Q�[���� )Xq����I���5��1k�����U�������H��wY�
ꝩ,K����|7D�*N�Yj`��~�-a����ٓs���"�:V늓Բ+�,3�0�t\�+I��T/gZ]�+�n�̖��h�M���-vE}��>���U�� �x5�p�%�	��͚W�,�n�5ʩ:}�UA��l3�iCkB�g=� �.7�P����Rv�Ns�,�M�.y�zJ���!�{ǿ�h�RrlS�u��h��I:�������-��� �s��m҂�n�z=�a���atE5u�r��e��!Õ��g� jv�Y�`���4!w�#�Qu�7���ϸ������*󨕡�|�8�|�Ր��5��"��`��9�m񞞄4��k�l�z�ͮ��ۡt,����	�� ο��� 5iɿ���D���f��B���1�_��61x��$I�r�p�\�S��i��I�b�2VZ_8^��[�c�?L�⯒�w+���|�9��O+�@����LT���e�}M�!3?c�bpi^ع�t	��k��]	%��Z�}�͖�s.D�]J���)��,[�����- ���׮mX��L*��`C�wIĕ��k<��ń����Uyo�zN�Z�ؚ���p5qHS��`��E�F�K��.������~���`��t���N��	��;Cik��,߻����V�'��o��g��x\@믣�[V&��c�ؓMc��no�I#}owPgC\��a���Y��G�K����6���E�p�^=}^�X�t��x�r=��yk?ۄ����p"�-c���w�W
Q��Y!��1�Cy[ЯdI�hٻ>�(ϖ�&|�����y�����0�4�I˕l&��63��>��V�NX������|�������[#H�ٻ�H\'G�%���𚚆Q�;=h�G��x��Al�?�M�^B!�d�5�눐=6��T�S�r{��~Uvv�k4�u�F�x���ub���$�����F���S����t<�~R��lTr.0B�H�}�8,���CS�,�4���T/fdl����ҲN�=<o��TY:� a]]�������ؗHDxMvR�֢�[�싉v���q�����������u1��E��#��ǟ�mB�/�������Q��7l%)�S3#/�)J�E"fP#G\�sKpȵ���c_s�obH=�ʻ��{�M"~���]��Q��%g{��?���@��d|թ�=��q�8����Ji�Iu獰+]vμJ4�w���� Ei�߂�-�g�_3�G�z�n-S��ޝ�!}i�"�{pK.s<h�w��"$G3�!�Mf.V1�X��3����!3ʾ��Q������F��*��-��Z��n�|�Xix�[�4�I�ؑaC�N�^�'�uW�~"���9���m�%���P
i�b{��9H�#b�y�*} % F�@j��!'�VAu�j�)T�'S��QYK��/&z�7��vܺ�B��[G��VQ����񉐉�e7,|#')���˙��B��#�t/$��-�o�~�.�|�%^����{���j�}Y^�P�o��H���%I�B���h���t�{����K�����>����g���tk��q� ���kqI�ę��͜oVzP՚u�HT�4% g�f!���ʝ|D\G|�"�v @v�I�H�X�@_�dk)^�M�ʾ�H�ez�3��֍6�,ۗq�4�'Ӑ�����D�����o�{�KV��OC����tS��4f�)�%�d�y���@$2� ������?�q �a���{�H��� t�Z{h�-?����ӷ֚7����C��j�B�Ht��REM%�aS����]�ѥ(�
��u\I�����= +7��Rp��[�VW����=�-�3�_��yyX �	�,C���4����W9ʄ��!:)�H�~�(Pr̦��*�ͪ6 Bl��?,&�ZQW��`nqN�<�Q���t"���F�({/��#l��>�;THʠh+R�������lS��[�!5�sq�I�"�/��h<��y^Z4g"�o�!{���J�ބ�zAϡ-?���֥0�w���W���Kj\@��~⫪.ϥ��H�qk�;]�O
z�Cq�L}���۸�'u�tP��ı`�u����x`Aa���:���oɅ�D��'�|殒@���Ե��߮S��k �]��E��&�~�?g���Y&Q��5���R�P9G�V��������:0�PRK���W p�m�����D�i��;����j��#��t)!�0k�ȃ�@{_*����"�ib���ٵ*M�*a��<����I������U�E�� 5Ny��w�|���F����O�:o��4`�3�A}G	�rv���9?>�.�XS�<���!cvD �
J��uhs)�X�ue.�pu�&�1����K.'��=�\d�Y�5���]m̠�D*y֥�%��@��66�$�zֻ�0] <�L�wnPC20Ċ�1`��wV0��u�
K.(�^[#
ȿ�C�+5�&a �6�����:����+b�Y�
��}KpQ+���Q��3���������~O��a�\�hMBiB啫s1�w*��7�S���D���-t�w����{vN8@)�)�F�\i�����ɕ�+&��a�m�R����h��H
����L�K�- i�+��W��^.Ζ}���#W�IūX�a����F����Tͪ�᠘�D�_?yG�!0R�h���5�.k�[a���s�Ќ7 JM���;���'���y�O�]��x%4���Ǘ>
�>���{��&zb�TT�
n{��x�c�0`���(b��D3��	V�gw�Z*�Q(�I��ho�	�L�7����U�H���X:�|�X�Y9�j�b��,�S��������{Y��:�� qG�e`�7�W�cw0@
p˚���7�k���&y��;q��S��ʮCt�I]�.[�B���Pw�V�}o9�.
���mO�_"��?'?�ʐ�6םҹL�Z7���뭴��U1l���"`�����N�Xa��� �b��+,�^~�d��vG֚�j��e�#;��8��}��^x����3\rW�0�,���KJ�)��b�uɊ�U�����\�%�D:��F�uj��w�&@���6]D�F�.�?�Q�������j#-x`��.��]B��A��7���%�	�J�սsߤ$Xo�'��<��k�q��P:�׈�I�gp��$�� dj�����)�h;��H��S�����* �����InŶ_��:�ws!det�,!�~������mӼ��p��8�8	��j���I��L3�	Ɠ�V�h5�O���~�F��^%ׇͭU��9.l�e�	�j������q|�j=�G(�O7("��J���	�;��_�<�b���-éTY�Qf.ф6���j>R����L>��T�U�����J���!𲮭G�|K�)B���"��
M:� U���I�XO��~��W�/{R8�k�.�bAo�WݭzJ֡k�v��o��V62�4[��(�	!W
#�yPy�Ո��;��򳶻�L����V���ݯ6��!����{�z�/�Z����M1 �� �l$�Ct��g��]F���ܣ:�rڕb�����4�pe�1)����׳�ّq,/�ǿm��q����p'�f���U�-Cd�i�x�p���'$�ϐ��M���
� ����C�v'ѱ1�)hU�MȒc�Qs��L�lD���͹'"����Z�Q7��>�CY�S�[�����=_j�R�E��0X����#�.X����\�o]����Gy�o�m�"�ɒoh�o�{f��DA��V���H�/���sZA��2��Jj�_%�Zo˽�a�c���OXY��+��ؾ�D��U����M����OL�b���,��RU�"m9��g�墂F�5V�ι��i��j��U&+��Хm��x���NE
�8En#��g��N��b�Ә�H��?��+g5|=!)U�s�R4}c80�g��G�d�����r��[u��`������x���_�k��3;�6���P*F��J��3��Q�k��S��b�1� bO\(`�,�w���re+N'�J8�̉��_<�ee�8B�e�4�� ?hȂ��7��"O�Z��<􁎒�G��3�_�ڶ8�ɡ�'���J����NT]���6��	`ƒ��p.b_�WԱ���m.������t~�&��ǿ]�_��[Ǫm�e�B�ee�wF��'v<�v�~=�f�0Ob�?��,GC�*�*Z�(&�CO_��5��U_d6�W"9��E�+,��4?=ؓ�D�����cT�P~]�ޘ�S'���Bn�;3�O��y����Y�x-��b���,���Gt]B�c��'88}�T�z�W�5>�Je��w�yqL�z��k�W�%V�D��wY^���8��cm��F�l�I�&��cY���~� w<�]�{gص�}n&~�Y_S,'����g(=�ި����)���>M��Xa6���;ANu�;�E@���AKV[��Nj<@4��� ���m:�����P�p�~V'q~+
��z�L�7�)	=��U�v�%=^�VY�{�b����nڡj�/]̭4ړ���y|[om�l1<���@�-}��`}<ƁZ�HԐ.���P����������Ș ���4�ؐ�%b��ߧC+�IC9������T�G({���!�J���Q�iR0��UV�
��/ �@�� =E�ꉦ 	�� x�5#:�0����,���Db5�'U%i���Rzm�]1�[�ܙ�V�À�-�:�V�F���7f�=�����x'���`�?�$�Q���э"� a�$e��%�D5�a1�?@])�����Ż���a	��O��b$�g��f���{K��h :%��고���^#)T�yp���R�����'���t9aۦ)U?Q��+��k��Kƨ7�9Y&��ӂI��A�79��vϔS!BXcm7-!
����r�!����>7�p1~(+��N�`��h�^�����ۢ|~��d�V|cDaH���s=����_T����O������C�m��èU�h@��:~����o�t�5���F|E���泿*Fo܍���Z���;�U�+2�I�4�B�*�j�d��^�L1�ёE���/}���憠I�5iC������Ϊ֐�D�(����x�a���,�@$�g�g���	��!b�Hw�yV ���PRk�8/���5��]�h��߄���T���c���OQ�1B�`�i��8��㙬{0'%X
(���(5j�Y<l��╘9���D(�>n�V�{h��y��/�	G1�$!�
��ҟJ�9��<�X:��½�'���B�G ��<��dߦ�ma*��a�����s.j��p(���7/m�)K���>���8;��Su�M_ᗲ��愝���	d���z�TA�ۂ�ɝ�F��^���/f�~���=���Ƌ�X�'�rX�YK���A^�����4� �#䏻d݊�>��O�e=�Bw�X�,�O�N��b+���lǥ��O\J�.*��J�>]։M
K���U'���0�@�CQ�i=0������X��r��1>�׏�����Asz��LAo�s��$37���;�3�G��om���"�1�$Kq^�ǔ��eU�l��R5P�u���p�Ҟ?��y�'G��G���3�I���'a�s�ZƖ#l9p���(R�U��w�s�"V}�q�Hk&K?>>��X����a)}j�]|%e����QS����'���e�J�+��qYJ|M��{��4�ԙC���Q %Z�˶q�7a`u�F
b;�R�q�e�ѫq��l����iF�
���G�~s.��c�گ#r����gK��_��+W��W�}�a̿�Y!�̖�%�&�Ԋ�#G���}OZ���- ����r�,����)��U�h�ބ��ѷ��
����dC��$�I��~f#�^�_�O�(�����'�BE2Eʢ�#M@�w�+��+W<��$u�ݧ�r$�qE�+'p���\uT[o$�e3�Ӓ�/�4x*��	�}HNU�EH7���K�����C ^Ptb3�Z�P�s~[�d���j���k�'�M�Ţ�9�,�E��n�����%�ZZ����]��.�E�X�/��S1�]��y��A�O����Yx�Q#bX���7S�"2�X]>(�8�=V�8�9"�0`a�f���@�45���C�&��ODk�b�����Ҭ�X��&�~:�ޮہP�P^l�h�o1Л�W��םޒ����:�p ��N�Ȓ*nT�n�(��d�h�[<H�\x��$:������W��W��j������xc����A�v�<����l���T��.����Z��"��}�9��1��US����דA�U�$�J9~n���\ٳ��I{q���<O�n��N�蟩w�acG��U�q��#�SaO�P�.�I��n��p�-�OM�o���(,g�%�S�X�2�{��NȊ�r�.�~��Y���݇g�m*��C�N>���0`��򖆋�0��v�F�c�:���j�Io��vn�EK����D�2^�h�g���R'	"x^��6I��3zR�NqC`%"I�N�\*���<�IɆ5&p�f����< P�e����=9�/��bL�����;K�`��y h7<�L��w3���3�dp�́h�D&�j��_r������f�Y�Z��_ѡ7��K?�((�e6�q�������#�������G������R�D);Wb�%	��.�%dRS�����������4���qD�˶H�̄�v�� ��f��� o�w��)�C�W���$����Wն@U���8�]t/��VÔ`6�stE�?�����X���\h��h�4C���q�����k�����/�-��OAy�ܯ���DVP��Ʉ�6��7+�tv��o�x*s��͕��Z�7�F�f����� e�n��� pq�àj/�N޽ �n5�ZWʛ�Ë�GJ�-�X�!ڈ���*�W��p�g˼Z�bs��S�Fl�.IO4p{���A�����r6�0�褠��@�4|ـ�E+Y0�ͯ_*ωq��r����&�˩�%v��u�$@���W��Y1KQ����C�J�6A�>ea0���h9�t<���)�Ȥ���9�X�Q���!��D�Z����Ĺ�j#o>Y��ln"wpCk�p�r<4�P�"x�	p��7��-����m6]s�%�[�!cs�9�s���1t�����Ia���9j��斀���ٞ{�E�	��p�x��\o��(��&NZq�ܻ�+.���
�S�9�U�7�,�P�:	 DZx�ݠ�6\-.e�FӚ��d�H+b��m�k�)��_�Y����Q,��j�'sLK���4��֌���l<O�Ǿ��*�$X/�$�"7x�DJ���L|zf���]A�TK�X���ﶧ��@����4F��v��/��@�k�D#̥�+3�_'�Y1t��?5��S�P�;b=�.cr@]mo���?I�N�Ҽ���Q��|��k�q�����\UL�̭��[�z68vc0�絸�	�l�?��`Oc��`4b-��(�|�����u�"��Q�� �# OR��$�"������]�ă����G�:�d������l����k����"v�&D��,c��(�CC@�D���OrS���9�H*8� �2��u���7ъvD�jP&��ޓG�����ȭ X	\~�����P�����%jՁb�C����jG��[�}�V�5
O��x��G��W���^Eސ
2�5ތ�Н�[\ Um���u��b�O��R�_������"���8ƾ����F�ˮ�4	υ��F髞)6�S��w�30����W>"�k�1)��������f9��#+�x�=/��ךI�=O��X�{�U_X����x�Y�s�/9�HV�x�~Z7~t�K�p>$����ӫ'˲��w4���\�\{%c;BɵXg�Z/���ϫB���?z�}�:}��.A�������F������{�8��c��.�SE\�r'�o6���(:��y{�ό=�np�jR����) ����t��e0�2�S��kĹ��3����LI��k�
ݓ��K;���/�7�Ã���O�na]M��E6�*���j�h~�6w8����	�Y4OA�\�l�J�vm�[������hDX�PQ�m���P�P|,���U9�Y�r���,>y]�J�Dl�T :(=�rKe��a��/.��];�����S=��T/�q!-i� LQ��#��N���R�vĸCJ��m����W�疖w�u�O��#e	E�jF�8�^��$�`墬`�-5�.���e�\�e���ha-�"��3�LF�[���\ݩ�&�˼����[�x)A�hNB��g���tT@>����y[EZW�̎�E�U�?ۊ���0�0L����Z�6:� ���R�oΌ�A����'~, ��
�����J�z��Uڢ �`A�"�gQ"�ܝsf)��6��S�k�Q��W��W#Fv�O�� �OO�<���rE,hG 7��w��`�� �X>��K��*I@9z4�c��u8�d. YV(�;�^� w�`�S�*h�ď����R`��-4�Ea"���`��l���
�� �i9�\/J	���vq�5�꼿�Q�!�����w@>yO�=��(򠡘�^�i^�m�:����RC,6��^��Ij��'3-H�4hE��H��G(8�m���i2o��Q�;"�TW� 9����T�����D��Q�u*۳���� ��.�4� A���w{5�i��],!����ރ�G;��q>��\�W��� �X�1���}?U�cbK~�L$��;=�X��ԾX�%qN`%����Egi�Z�t�}����W^A|�$1�3=#;	Ukw]���t����O�f6=$uJp٩)�k��3�Y�zU��^ByY=1��a��̖ةƂm����SݍӍ�I�_�<3�PY�,���6�I�F�#��ic�Qչ���J�%�@V?5�n��Ջ��*��p`���a��]W|3��"�\��ch�R���E��Q����2��T�g���6�)@ECw�n���$��'�S��a)Ύ�/Y8~_�2�?x��n_�ݎ���19`��O�4�}�7��f��6������^8NO +f,�
�@>�������Zp('~�bx)���(KJ�n�j�-�
N�<�%öp�b���̱J��/�n 0��Ko[��Z�9[���I��򵬋12񔘒n�=�"���dy���8`�N:�1�U���rNG5$��~H��,χw��ƃ��+?�U������Lpo���PD�����HL�o����!��F�,X���DD;�Eq5����Q���S���ъ��a�ݑ�ֻ�:�t� ��!��Gy7��������_	
D&�f�<E(lx�R`W-���*� �#��po;鶫��=)S�H���񏒘b�Ɓ��6ȃ��l�`_b�1�^���,d��DVh��y����n�ƚ?	�;pRJ��)$s�&���M���*������u�s�U���� �5T-���f�������=�Lؽ�_��E�z�-��d��W"��Е��5a�p�����'�T��tΒ��b�`t;��*����9ft�^�"�p=RA3�-��41`�yV���1��۪=�"s~ӎY����I����ϴ�sy���` �(�	�D-ׇ��zg�t���.1G��$��젶���Pۡ����:��/ܼ�E�?��q�B���� �Vw��i���>Rr�@��0�>���v22��4�$�����l��-\U��N��;����-�W��OCͳj��T�M�$�&�&Mr�/�")ݽ����a��M񴲯�A#��������~Q!�K=��R�́�G�
��d]��w��x1�E5�x<�2J~F�%��mk7���j�/��F��ʒ!�}v�e=����A��e����'�D�.p׬��1��C�]�y-vRs�K��7�@",�"��ut�2�!�w�� ���
��:!něO[�S+����@�yUAA~�ϭoM�e{5�\F�z)аzv���6��L�ܐ�JÛ����
�� =Òn��]i�C#O����ɝ�m��ML��k@떇&�=�M��1�ؿd�;�˹uwG�d�M��M0�H�?L܊06/D�L:(��8�v��߯�j�_�"�(�+�f:a4��3���){\�h0χ:���|;;�z�|�l��MW�0�ZCӫ}�h�|��,���M-r�#OD���aީ��*6Λ���Ԃo��ɫ����W�f2�zŪ&�h!�a��V��a��P�'����3�ϊT��h�掊5�6�-RX$�+�o<�$��q�ov�΅;���^��i�?}�V�g>/.��ilX����M�,(ⅹk"�c]�ǆ�7w��Ea~�D�`��6�l��FjMW���H>����ui}�XS8UNN��y�Z�N�ϭd$� qH���X���OLRT��/&[����6)�
���UD�l���爰��S�~���ױO�����/G�-�2煛�?!o�v	d�� j��6�ѩ��s.)��X"��<,/'�Sm�*Y*!֮/#T����݄N�L8�@CЊ�-��*jo�<V����r�z���}.J�MĢ\�0��|r
�������Pf��ǧJ��VVɄ��D0��w��xP�t�j*�#��A��&݆�L (�OFh�o���\kuv@�]�E�ڮRzS�:���	݉�E g>i�6?|�����Y-�+J*2����E+'�uc����� kZ35�J��z-�4lj鼐h�β(G��f��7��_Z��r��>����F�3�0A󎟡��Z���W�Iy�Z�L�R�y����r(7B���a	�s���s�Zy� l��������
���u��3��a�l�a��|��ں͏�3ZGo|+��Vϩ�\/;���V �b0�o9�鲌#ױTҍ�+!:���FͰu���~e�# ���r��������?��R�-��ƵFM�<|l�p��i�~?�a''�,U�0��瞟@�&!:פnϜ�8z��)ڪ :��ck5�kL��H�LkK�f��`]*1;/��a�W�+�^N�xe_#���[�D�ݦ��k��8( ��wn=V�g��i�Q$^���ppݥ�ӼidE]�3����%�,#*����c������w�� u1mq���m��܃Q���qN�᳭����a���U4q@�6��|���Y��E	�W�J��t���� � ��?�����b&thܫї���v�9=�y�C�/��&��s@_�X��~�R�'�D������3m	F9[Ȗ�h�/�рx�N��s���|��ͺ<��p�� O�|�#C��ġM�&�l���:[B�T���	�@q@֤�a���o�O�X_���E���e��~���W���;%=ah2��;p�g�l|o.�c�E  aU�����LNpd�1�#�n��z��I�d������{#�Y��f�̋ʖR�l�aL��\�{�A�b����F�`�Q��q�#���+iJ���+��8/��+!�.eNu<UBSiF9�ȓ�@��ϸ;ދx�4�ri�fR����H�H�&K+Ci�n���ⱔȤJ�m:R����z��`�S�Md�;C�";�(3:��*I�R��'������o�J��,��;�"�J�RP{ڟ���
[>\R�R�z�A6	\�s�1Ý�M�D�&�n
+�|���S���_��t�y����<��J��؛��\O:6u��9=
�y�����ƍ��_������y̡���h�fq��tSS�;��A��FY���i�r	� Yt����K�:%���i4�9k#��������A.R�o@e&M u�,#��]B��W�ܿ�2���|n��Aۺ46Dv�{�2�݀� �%S�2��\�	���� XO�XNg��m���z��ފ�Khc�m㦴�Da�khR����]k�~�Q풰�����g�����9�6AǕ�Q����n�|iDEOU����no����1��1��^~��	()�_�C�K��5�U{�����DϷ����\u�}�%��A���܎>�SבR^<����l��kIH��M��$'��h�����` �о@����C��U7��R-D��?�M����W�~���yCy�R2��@]���Ё|?��Ã^q�K�˦�3�) �eC�C�/������o%��Z�Ψ�8fC��H����a��91�F�0�o��v�@�Ӯ`�$�1_������ �]��q���
�Cֆ~�����v*���%�p)���k��Q� 	�����`�Z�*��,�*?�\�Ǭ��v�EQAJ��W >5�4���|6
NV]�l}C�EC�.?��R���L-�w������I��7���C=���k�h�c��#��d#c�fTC�E	���ȑN�n��2��s�M�E���]'���Z���H�v>��gk��$�X�|��(����&����BJ��<+v'�ީzp�䖵tP�ڻ��7���j�9fcUc�!�۳��s�w����ĳG2@-�gi���@b%!�D�k�{qEJs�?W�h���k���q �5��������s ݏkJWF�k�6���R/4���)'5}C&�|���������tv�&N���G�jG�̅{U�ܢxb��>v���?/���DY��!9'e�R,�`L6��W�W�Z�������%c�W�Z��Shc��'�{�ת�[2�ʺwK��O��J��)�
��I4�����)��4#V� ��(`Tw�Uҝz|�;�%����oō��@���KI'�H}*��C�̮w�O+焎�� �Wu<�[t�瞜��`��΋�m{���\o�]�޻�����BJ�A�r� �9yF�wف�1���Q5�����W�%�}�NmQ~U{(�
��J^����DSw�1�y_' �'�OVL{�14_w����UX~������������@�P@��x���(�xX�����"�j�[7F�}�`Ⳮ����y�tݲC���AK�g���u�y��ey��+�>]A$E���B���%}�dM�|����&������k���ujc��w�D��l�C\f)Wʢ���y����4�2��Õݼ�w͓=��1A�{�tL`r�Qs˥~�jR������+s[�c�<��x�x�"�F'��}�0}�O���IzjX��*�(� 8}�2��n�x�����U��FgR���)9���e{D�u����#�!1��e�h����ӠE��ďs��`�τ�60c&s3B���5@6�W�IX��Y�c�����T����� kcDu\ ��3����E݃�5�D�k��)�"|B�㑾��U����S`s7��'R��wV�L X/2K�-ш�"� wR�����?�i�d맋t;b���ŗ�.\�lfax�	;?NטD>&��K��!�E�I�����9���nEQ��UV�c�q	�n>+2.���O��ףC��W�U!�֠�����>��!~�/��6>mמjT��.c]o�G���!�����g\�*4ר�;7-}����	dh��@M��hg
fV,ْ\-�'� �� �j��l*�C��a��B"%e�z	*B+���A"B����s�=Q�f�ј+V��������(9���R׾�6�-:l���4-r>P�Ҵsa�/�x�������FJ�B���CKZ�83�ifU��i�Ϸщӳ4�����Zm�
���c���M�o.MK.���85̱#�d{��|X�H��|0q�6d�37f6�3G����Z(n�H����L.���*�]�k�=��nD$�}w".`���z�YS�9�2Ƞ�=�������n��~"��ї�;��?~�����5�d� �<��tpwn���bӤ�R+\�H����df�,]jVU���va���	N׬$vq�@�$�FxK�EQ�cxZ�U�S�9�\˧d1�To�]�aj	�T�BN���M���'4�o8�o�0p�P�[6���g��&N����ձ=�u�;�x�E1�mA���2"#!;�����������iWѼa��Zla~X����*w[�d�$p��� ���U�ۜE�]�G�\��Bb�ɬ"��v�	�+���q~�|����Đ��a������A�?��a��G:f��4'T]>�%���뎎8#-�#�1/ޱ_[������}xb������2o%s����v�9�B@�}�F݌�	K��:T�&JP�AJՔ�(����J_��%���,�w���A[���+Jb��<|�[=I�h�q�@vV�|��@�:��n���w����C@��0%��b�Hb꼴�_}l�%`�e���36FFcl�/Y��v��O�zyIo��o�X���0��,�7FM
 Əh�����R��Ƭbf<س��xɱ���4lg����`v�zp��ė�3�X��Ow�iU��}���N�먁�7q�/d�2����@��]�[W���󔋈�&'��mj��r�:���'�w�����x�����ne��N���5MJ!{�� �[�oG1i���j����۹�8�ز�_�m�8(��������+;��n����$�X�H��2Jw����>`�e����F��ǉa?�a$7���5,�Q��
�#!D�*��eT���y��@��`�����t�y$��=�2�+��Y*e����٧}C�H�ƌ���L�B�U-r�;�
�z�����Ns���P��>v����YnF]�1�B^�e��7�u������7�R���.��B�v.��z���p(qG{���+��Nj��`Rσe��e�_�)�
f��JC�]N�������jz͢n�]�2�����k��3B��x��6'r��aFݤ33��[0��)��/��V��k@�����[i]�� �P������I`)�)~�ީ���������bn�}D:�g�=���H�i���퀷�d�ndgU�_jb�;4�פ*N��?���1Ԁ�@iG,�:A�6���/��K�.5-	�ґ��#����,��}{������
��1<�!.~JO�h�b_�Z��+<�93N;��W�t[H��J�����4����LO�h2pp��;򺍰��i��ܟKH���ܸN����9����c�c8�w@���Q-��v��r	V�H|�ʘ0��N����M���@.�](#.�+璱)�c��S@��xi!���`_�3��r�J�>�fS���H;dVt�к�!�YX�4�x1 8���q���x(��f����ϴ3:-Vσ�Ed�CTv�o��b�E��ς�3nQ:��<cq���H�%T�(��uk��{ؠ��T����8'����3��ssx<�tJ�!w��}5.���߳;��,=�m���"NO�b�i���V�������G>@7���Sͯ�1{"us�_Sx7unzbyW��b�i��t̛[&�*�+t�E$�O��n?���Fv�#��E\��{n}|D��1N2��N�SX��<V
���O�(�_L��&���~ =zX�m��ڧÖ��-�Ԕ����A���z�1�$f-�"1��R	��W��Z�[C�ra�p��,ǖ;Z��OJ�7\q��ғL_���5伝��YIa5�7r�J�B�s�E�і� 0&S�6��CQ��	���]����hs��Mv������h�*h�%R,��'M�I?��#�9[sǵ��3���X*�ku������;<�m�[Տ�ؓh�{�A+���b	t�]�°��kR+���1�m��.���<�v.�oH���#��T�
����ݐ����ܖ9*��4�����~���W�;@0�)�;����,�@.|��ϐ�S/tr��A�W9n��v*�"�3�t-c[���8���2�,���aܸMe�����k������K�Ǔ��
ܮ��U�4�م����0l�c�!-��JH�Weƾ=�3vu�S~�O��>l��8�����cS8;^�l�!/(?q���S"��`��Ǽ� \%�8^u��4�}�n��1���H1N�;'g�]��z��I�;]�50`�ݩY�� �W��+��9X����$�.Ш�����R,�/U����pG����I ���(?��R��'"5�W㪎Y�h?/��Ѫ�B�J�ʩЉ�PZ�r;�uێ��J&�j�u�F��$ +�î�́*4q_�#��XV0���>
���k�F�4��/̈�~W�I��l�)-�d���
/%��hWhf��iJ��k�����+�u�J�"ޖ"��Z���:a��s�<ۢe����Mv����a�h���n�}h�Zb[9��}ʅЩ��Ѡ�*Ⱥ�>��-ҍF�n-���D��-R�X9R�$.�]XvQ�9M��|��2��L�7��9�E^����㧢fG���s����I�w��$#�f���6���~�!ۻ0��c_#��{L/�:Z�1 I/��~4�F��c9�6o�m�o̚���"ι�,���ٌ*�j+\��X��H�r�O�[h�2r���<��X
���3�����������9��_��q�)��q?��sp3��·�0,p���f_ߙ69�/)�a����n��hd��������,�BF(�q��1곙�#�M��Z���'�7���,얾���}��o@�d@�B�&r{:�C"��wB@>l(wu?��S[:ge#���HÞ������c �P�u/�<�i�����r:���d��ON8�V�m3�9��7xw�?�'n��qþ�Q�,�B�?�� ��p�^�g��A�ǽE��l6�>��׬G	�4Y� e�Խs�8�c�lqe�O� y�,��HV��U�i����ޅ{��3�' ����ފcJ�_\O�wrU;�&*��u�d�ɗ.�a��;��j��|gf�xʦ# ���QG �z�rM��	=JZ�`�t������΋�B�.+G:�am3�����>�b.���!6Gh�<��i�t?�=��v�d��؇hng��Lfo=�A�a� �M̺���G%!;A�� �(�`>��Ͱ�`��a�ҷD�:~$֌U�p��n���S����\�MU	�=k�����J�AUO��$٭�G\��G�:�#=d����9�����ꪨ�f�c���{n9�k۟�ĳ��6Z�pt��9�FN�~�{�r���T� ��\U�F�2Q�v��1%PƟ�͐�4oN�y������h�9,#�*�}@d�� �y�m���1�+ ��IT�7���_jqڊ�0��J��xa��h�%m�?�쫮���������c����q䤬�ӠϽ�ZecgK7`��aF��Ȑ_қ��E�e�d�Pڳ�ߞ)�<
��5��V����}��"��cm�>�!�Am�x�I^�#��|-�N �@�&ʤ��o�×s�EZ,h�������=`ud���Z?~�o��#�1��V�!�En�x+E�Ù�lt�
m;5;��kS�Y��Jg7t A_���
��t��aK�;I͒�zG8�[e�n�<��Z[�t�6q0�����c���.�e/-#���+V�R`W$��t��º_��r���^"ↂ充�'ܓT�mw0�n`X^��4�S�=�?w�w)��R*�H#a��{ ��t2����񋠓U���ê�9�9X��)J�e���EɎ3�.�a'�3��b����y��&�(F�I!1�������u�iW�̚r���,H`�'x��*�bqW��Ji~�5�;�>���-���9=��lw��D!34;u�)c��U���*]�bt��<��ӵwN ,�CS�uW��'�GJ���6Q�����N��-������	��+G�%����{h6�xjh洃w�[w1wq6� �����LW]��7��V�qy\=��+��0�:u�d`�
ʜ��WS*((&���)>&t�	�ٯ�C]�]��k�d �}�U�8���O�kxS>�i�{ҿ"��ˁ�ԺH�œ�M�~��F����vB�I��]v�?�{����E�(!�nnM2��lE�y�*��+��3N5Ə�@5�IF�חb��0]��.����R(��������*�YU�� !�绯��ϵ\�@cc��Ǜ��"2���|���(�$NP�3�2%��kjb �d��wH��Z�,�*DԊC���E���J�?P-�s7&�'��<��u��z��3!��G�xw�>��tnJ�XQ��x�5�@z{�������:����:����}��b�q��{�u�
Mj��]{+�@Y����S��oJ�]�u����d���+����]Ab;«��W�F�!���|x��i�'�3j��U����-vd�%�4bD�DV�I����+N/d#�r5;"o�.���e�8�T�D*�S��O_�sţ�bG��������֧nb͠/��&�!�&l*�*���e?��&X��/*[�:�_� ��J�I/\��jX�PZ�DL�8��͵<�7�5N�K���h�~�=]���$�*������nO� )TB"�3�y�Z!
�q�ջ���A��b�,y)H�㖩�Di3�� 2���<�Ʀy�uh`K����f���|����~�3I*�N�+,�05�P�����:�VY�������c�

�o��m'6��G��Bc�������Ҡ�hh9�@ٹ�G�`ѝ����sQ�P���ţރ1�Mr��R�6u����0���m��*tј��K0`A�	�r��dU���W� y
w���q�<͢�,N�u3 �!���`��?z4,5Ymi7r'�DC,���̓&�.&o�H�
���b,�R+�0dEH��_	"33cDOer����y���P{�b7Cx�\���DX�O
P;�k�G� 	
`�	<0���н�Cl\���ۜ��.���q����f/���^����4�t%o;Қ>�U5�3i�4W-���b������N����q�\�(?��(�S쓅8ܷn�IA�Κ���r|J���b��駁$n>+�g]�����U�*�� ���Itk!)�&f�ghV��XKM�6�ܤP�`�'yW�L�����.�W-���<�ZIz��P���A;�"1�e�YfY t#{Eٓ��c�L�����m�owe�Eh�l��"f�ƹ1ۻ���@�:����=�am�1̿��ߪ��w�6�%V��"1�.!�t��㏴�ON};�	��&����ڦ��ww����!ϕOPXb-o�`�t7�,�E�����W"�y�2��ׁ�Cї}J����Ɲ^��<~<�����p��P�H̑EW��r� �`�Dy�sI����6�����K��!�\r�h.�P��j�R���h�����)�#M�1�M9A�\��mG}�����=l�}�H�can�AH�?��&1���v,c2�5݅s3;��{��7@�p2��,JV�C�c���E`0��g����Y���rj�vY�n�I�����kw��� 4�����[X�&�Z��w�#u��=D� �Iy�D�3�ӟw�z��V�����\/�Ӵ~�*����D uq���:��ͳW���<��Gm�`b@�����̥�s3峝(�=���c2�>%RF�K���c)��k_���"24�s"(Aj!F !����&��\���IW�ÐܵuQ�Ea�|\��4�JW�����7����UZ��@Q	����Y�!�]��^���q�ₒZ��B�į��k�����0t�qL����p��|�^7�U��7��_)[`T��5�-�*:�v�o �~�L�C����]��X�ʨ�@������b�*��'b��ͽ �|蘾m~"@��h��@���l�&�u��K��N�+%4���C ��G�?����V,��]�Y4޵��?9����Pu�ۑ��g��`������Ԙ�%}����o�hك�Q�u��;E��
}�
90�p�Y��ʉ�/]XɎǽ��K��t �}�������Óږ)W�����ҟ��:3�����8۩1wN2��5  �\��n��i >݀���e�{i��#f�;ߙ�r���q>�Ǹ�l��|�R��mAu��w���&Y@IE��C7ۣ�'كjmj�����������Q����*DB��@*>Y�X�x^��.��uC���U�b�lIJ��
��Hԝ��dô
�S�Ŵs�x �h���C�=	�v5�pp�ii$�s�U�iO=����A ���*%��ϥ��{�2jO�	4tn��d3p�?6]հ���3�{�S�"O �
�!�L�<�+�o��rb����r$�'�(�8�v��
M�(�e�=,ֈM~͘�}����5{�<[���c���d�ђ���f(�x��o����,�P�Ř��e�5ܷ����[��z��4J,��l9X�N�����#5\��Z�$�~H��u8�&�8��!�����߅a��~�jh��ìB(P� T�/�DV��/� a�|��;�6~M�R�{D�į�Ξ�Ё��5��0!�v��3ou;8b�N��@}l���
�`�r�#kTp�f~/�u�kEH~@�]�nF�j��ɧi�q"��eC�Q�p<��R ("��Bx���X�H&V�^�;F��y`+���c���/�Ws��&
e�&$��-O�J#OS�p��R��o6L%�|��+ۗ�ϰ�]5nv�k�(�^w�t����:�
� d�6��6���HS��gA]~z6��U�G�Ôg\Zn"������{^�d�=o�JI6E�.�r�F��%ţ���hϧ$���3|��fb����S����Q/NE�����m��>g�
kFW:O*�P����{+��-����i��m��A������z
��@����t��9-Ț��3/^��1jP��3`�p����YH�_�n��Q�?�>�v���di�%@����\�7�G��r�����}��U:'����)0# I&wj[���l�����
�����[,���'���k����~������i6A==��i�����W��4�H)O�r*�F�	(�2-奩u���4"6C׎t���O�D����#�eFO����KK\4(A�*�t�K@��޳�U����#�MMh�~�Z�իd��wN��Ǹ�u��z���Zs~'*��
�d���HB=T{3�(�t{�%�b-��,�Bh��fU�`�!�!��#��]e�f���CP����K��Z���c��6m����<�{_�@F{y��hM��чr�mU��'N����;��S��5�yV�d�M�:�m��B�-�R6����1�
�;�jF��}�7���6�a>�F_�'>����zMb٨y�X�=��d���Z��n�g;��A���Ν�^�+m��Ty�iI"&c���/I�N��[\�bu��#2�Px
��	��T�W!�N�&=��3O�ab{e4�F�d�0�[I���>���8$��-`'7�rwo\����*�2��c�&#vNԒ�6S];��Wps�߽y�(���Ɛ8��)�!�p��3{YW�C�d�n숩��E}��b�� �:�/֑V��c��/X�(x�W�Ɂ���� �I�p�!�,�T����vݳ�.P�I����7�����n��R朚���w��������$	91�Ǵ_�o!���.�~zذՂ� ��w��`p����!�6��5�4�Y�}ռ�)+���m�*eu�h� 3�l������P�c�����T�@T��V�<tn��+����U �'���&�� |y�V��0:����1�Yu��K��/�\m��s\orr�j�R����;��N/#��تk���]g�n�31>N�!d/\9��z�
��z*�\(�禞�j�Ȗ�H��MK��w:3`8��U��ub��ũ=���S���P�WA�s�H��UDl�/Gt�X�s%l�J�U��=�����Y�8���7�yB�_��Y�SM��{Q�A�|�*��0w�U��=ĢZ�~����cl�aW��Җo�H6��/gQ��%H�:��.�����ɨ�� �����<���?��E����rUF�ҝ�`�D�Ń��Ԩ.�f�v���pwC����Q)��G�P���/k�gA��������7�Z��Q>�ZdNc�����f��Ŗ���=6*��QT�A�4����|Y��XR�)G��ތ
Ȕ��Tn�k*���� ���2h�/�f��T������ϸ�a,�-LT4���C�6a+|���텏N�ѐU��e��������&ҙ�t���B�L�6.Z�L�� ��lN���|:��X��X�
`�j�h�[���m��M�awOװY	o4��4���!��3������)�bC5�
P��#ҩLx|��=�۫
Q���� 5�-���]`Ei��
���6͏
<+�@�=���]��V~�]��7�P��0X��zŪ���e�G�0V�fM��bD2|�3$�����{��ףԮ��^J4q0v�V��g�ju�q��׹-k�Y�� e�&HP���a�똿-��2U����%��Z��R����ꋍ��/��M�f�G�b�uYzC���{>_x�t��<�D����ѩ_����fWty-(o�ʹ�B ���	Jq�@]o W�_(��ĳ���2w5wF��"���~ᔃ<�mE����U��N����1h�b6in a{xn4�����	�������N	�nA} ���+oB�I�W!�'��^��(�hH�,=��Ӯ>���}�1s5Xr�+�֙�DD#�Xt��hA��M�t�	�K�T5%}s��~ͬm~?3@|	 ^gkn�҈�j�C5�V��<%�X��+�<�|����4�ѳ���cXl(�X��/��.�Ek0��;�cvK�a����A���qC�2�ˏV�=aPH>c=��f�8�2�|��5�f�Y!�����	@�T�S�A7w�m�8x���o�S�+&F[�6#7i��4�n㙫��U9�0#ѠKM	~�K��rO/��D䩀ݘR�k�e�)j13��ݺ���Or��"��d+�n%�{�k�CR�/��6�'D��.UK�Ĥ@�c�H�}�%ˀK�?$6I��ԭ�����a8�N�S�}�����6���f'v�;&'5�d^�<*��f���;[��8^P.�ÕD#���\��2k��@z�h'H%�1���r�_��y^ݒ+����U1���c}��M}��"���S�3���q���?E�S�d�e�X�ݷԻ\�s̆g ��<�e���!�S��?T{ㄣ_4Ȭ�:�"����cL(ނљW����e��K���jKT��S�b�����Y��a��o&��fv7�����1N�tŚt�ʫlp9P�U%�?N��e.}�#�%jl�A��r�S@l��`�mhu��wn����TH�
>� oI���xr�]_�y�?��~Y3ِ${���B�+ۻy�"����3���ڼc#K�� bq���=���^��&6�~ō�7��9�0�55��R��r��Gvd���<�c�p͹I���Y�P����~b����P�{"��-�_j�� �������p��[g�.�1�V�JH�PS\����q0?�i�>�2��M��QǓ���ފ*�R{<Ui�>�	�0�x�?��/R�������U�jA�=+���Y�/���;��췝�<;=��@�`��mxl▎vx�O��:R���i�<Τ}5�9�AN�Ŭ�0�J��Il�Q�u[:�\��ğ8��L�%���*{$�B��v.��?�����LY�i������\��/L��F�����o�Μ�m�����L0v�GP&U�����-�GL��\�&cM)�#�7��
����NOڱ�&������|�����I#�
�ef�O@O�r�o����FJ����	"��-̸�(*���x�r���*���NWF�����uے��z/�c��`�gy�����?*=����aRTF��Y��'NVy6/��X���|��O�]t�$�������-��ʳ����7sfD�*	O������jBp_)��g=i-!���*gsl�Վ%��n s�o�yR��Gi�熝��m�|	�u|1ē��
N3'Ψ�x���k�Eݣqj��9�o�E�1����_����S=���y��E����Γ�[�o�d�u[�bk %���}�����EW���Kç/:m�pd[��Q�y.)�[�E_�i�9P���q��'nB��=p�6S��H�c\�ڲg�^Mо�:���������}&^��<[7	4ݝtb:"�t�b;#S�ʠ�7,�.$ƞ�~,��<x́|Q��h8E�۞rM�-�i�{̨0u��&�g�,@{7�Kۀ��O�x#v�P۪WV�"��O'{s��p�M$��n~(�������$�(ӓJ��6����S� N@?h���g���E�Lf}�+�:��L���c1�,p@���B0��y%|�RB}9o� k�K�8ܣO����*�b��'/O��u���=���z'�Y��|���s��r�]�?:@�$G|�,�'O�.u
}�z����w��@t�k�oD�s%Vbة�;Q�\��X������S�SU.���Ny��o$�P���1�&7Y7�	BP�2�*v8�
r����rqc��x�����bl ��ͪ�*��2�����(
����Q;�I��멇���ȤAj�A>L���j��z�&EJ����=ܜ@>�=��{�c�@P>^"F%�WN�$nk�r%%-Xk�����H���$u7���A�ܟ/���[ ,�Fĕ���h�\�}�'��(��3�̀�G�Q̌��1W��R�5�m\���!����D��r���s�QJH4�tf�WnL�DP�H��?_�jܳ6�Y�Μ�N�P�ger��Z�P���V�[�M�'�!d���T:K��o�ĺ!���ӂ@��\�;��9l�k��,�r~��З��Hz�nB�;gؤ b��f1�;~T�KH����� zH�hÎ�����ax�g�"�~Y�׃�T�R}z����vc��U �L�
"8�7��^�a1��F:�߷oއg��޹w���9g�^d#BD�!�G_�C�GG��`��C6��q��xAy˙`�����נ�O����ưȬ��GJ�b����/˼��>0Q�N����,��&�m�3J��,a�ˆT�TLzD�9SR{���ߍ.r�$+Q��5?��t��Q��{E3�|ߪu�y�RxtſGՅ������B��|0ޭ�9aJ����Y�~��8����ԩ�Ye� �f��3��_���?=��|�OIkK�/æ�{6��&V^ݿ�7�/���k��H���Lu������|iP>��.���K�t-L�G�8��M̬J�t�u~�׾��gq��\�S��SH�����'��`��7��S��1�r�Z�ҙ���z���,����t�csm��21gX�ݭ��&��m��r8F��Hթ�&G�08�YԂ��'lz�N�B���V-�y��%����RVZ���FX���=r�@�Cr��ei���Zݬ�JE7�ڎ�m|SmJ"35:�]C2j�8���j����cm�:򤃍y���-���X���Gf�b�m4̤e�4����zyK�����i=N׈̀>�������h�J�����7<.��u
�9�(JҽN;����� �P�a��;��n���z����N8~-���\��<?OF���c��#���I��,W�@�mz���j�qy?-?M�VZ�nK�/4{yRD�.;�<F�=�F�t�T-;���r��߫�~����F�0�h��K�o�xƙ��76�h�"�KNҺ4�zDߎf�PRrQ��(;]��$��x*��藕$�H��$�*� �UT����g�:�<ŝ�UG6Җ�k04|;K������Y�]KU���v֫~��}�[�H�h����Gm��A�|"C��Z�qJV��O���IN�W??{j�n�z����$���E;#j^2=��Z�ɾ���W��od�����0�B�s�އB%QR�X,u�}��d��b$_	X=�ܗآ��`�
cX���2:Xc�rkb{�k�$8����I�Q�c�7�6����ج%+,%��sJ�J�m��ZN:=�&�5���!�n|ꔫe捱N�%r)u�U兽����k�]�6����N2~�,��`qn*D�V�ދ��q�au<�� ">o}ڻw�b.��vvi'��E&);~��O]}U02�%�.� ��GO�B�0�[Ɍ���m� �9�	�X���Te=�)I��̌�x�D�jpt�Z�C�y�`�X�-a����D �!��l���M��dG�lZK�
��/�m_q$�g�=��jJ���$�"`�-�҇�VI+o"�|�N�������E�xȷ~��`�3�6"�2p{��
��"���ׂ6L9'׽��!�#?��� j�K�VTܣ����� S$J1PB�߹�e"�n>6�\}���v�@k�6���(��q|���zW������8��/GJ�����*+�v(^E�THM3��s�p�ߛ�vo~����Q&��e�{`;V�5�U�Zs��j-�׃�8�@"���L2���(-p�M_!w���
�J�K�jU�_���9TK�d�6�62���1��H�ܣL�&3T�܋M9N;�"�} 8%V��$�1ٟp�k%#�r)~s�F^�;f��^���O�7&���	ޮ��0�I�v�o���X�K\��oZ�2�b�f�AC�xDQ���r��%�N�����ʩ�.u�^I��5*���o٦�̝1&�{#��*�T
j��#f�P�U���}�2��I�6씎e�lH�½uW��w(�.8�g ����b���L��k����:�������d��\�3�x!)k�	6 MF�&QQ�\.o���$,������O�u����f���w�O� ��Q�TZ�Փ˲����RG��Bkvq)��0�nO�����O��v5$��@P�Z�E�GX� �(ߊ9��,S���e@��da~��g��"{�j�[�[|oFɈ;�Я�i����%[f�M�c�$���*!��5���AOy�.S|E�KP"An3�irb�п�-�#�!3	�V�����m����	�+p���mz�"^B��4)���<+�ܼ��v�w���n���VqD����z�+
c����}�NbH�� �yn�i_K��WU�Á� ۫�<,�D��]���e�\*�;"�����ŋ��o3��Ly7䩖������'�^�Gb�g�Q>��1?�LM�ĥ���GS֛I���e���A,��VA'�@�Mf(�x~������8��t�;�1�؟�A^��1_6B��p�[ȫ���M���M�S� ,����Nီvtnr������3����5e�W=�ˌ�D��$�gG��;�_�\��[z�,��+��ܗ��FM{�,cj~H ��F=^��B��[�0VcЄ���������<�h�ZL�2��<C�:V0M-����1v�OW��abgVw�Ő�Uh��G�Ņ��y�u�%���yX^_����n!Gk}�2��L8�x������ �Ǒ7�R0�I�JVٻ54�)�Q׌�@�J˃g�F�ey�B-���l�a���9̈����|w�h�s�Y}�� ��2Q	�h�S�U ۺ׈�XW}:&ŬYeX��z�/S�6���e�=UuG}��.��܋zh��HV�(�ŭv?�X�Jp�p�|B]���aw�bΑ}fG���שe�ζ!�c�j�U~�Hi�,�5��}����J��ܟݬ�����ݨͲgW��_X��NtZ��^�}������i�Ș���8����C�J���O�w�:
�(��D�0�.�M1੯g]P%��J����1 t���3�狚\F���W�h��1Әc6^C]�W��4�y/x�(���Ɯ��ֳs������$Yŧ��n)h��;��͢#\`9�K�. :��Q<}Џ"����B��1z�������ms"z2�1a��`���!%j��k�~r���8��}�*�޽ջ�|z̳��ߺ@]��Y�8'���ƞq^�>����σ���2�2��뼮�dyÏ۾[��7�m���Ylo���z�ܷ^�$G��41b�j/C��2[D��E�V�E��=�j�.���Ɂ��I�����놠�هp���ݢ��`{{-��8�Ԧ�����xf,��}q�OqM�*����`�DB�����J$�Ka��߇}`nΊ� �������� n�SrW�i��s9�h�J��UL��?�Ђ�x^��>�]�>Z� gߊ(Zd������o���晎6�Y�!I4��23j���&�g������8�Ӗ�gރ��a?�!u�ar��h��=������\U�>A9kll�!c��L!�p,n��_~���ɗ��U�X�7���I�����"O���.�R�����SOV��K5�a�wT���;T��V��a�1B����8`�$K���T���.�Ƒj����������Ӹ=,\�J��YD8���2Tp�������ictD��}[���Q۸y�9\�Y<C����]!O{�y�]���G���lS�����_�}m(����b=~A�ǽ>a-#���P�ii;��Sb�w�_����Jo�� i-c����_];P��N�/��Dz��bbՄ��X�W'7�������jdW���<|zP͐/(L#s(
5��.ل���'��t>f��aa��tSf{�=j�@�H��J����|(�59>GK��)����.�8耻G��5�]qN]O:�)� {$�g��N�M*KQ��������@�- ���fS+*_��Q�^�8�BZx��k�RcR�Bi�uU�i�5rM����ElB�Z�J+���S��7π���AB�v�� BQ�,F�v��:e# F��M����}ʄԐ
����]7k�c%������~9�B�c�x���ͻ�G������ )>�f%;Ys�`�&ٙ;m���?�R��X�Z�ڠ�}S��O0��h@9r
Ku¬&�4,��2˖)����:�q}��ѭm��W�����v�f�9)�(��+`#�V��ȅ�x�~����CZ1��	e@�uZ�N��!�Ԝ��U#]N������?m��=�_G�\'qIg{�Њ#�R�92��r%'>�Puˠ��L���|&Q'�,ŁHl>���z�R\�3��j�Q��vm�؈. K/���m_� 4o�굫$�"�j{&1g�O�N���G�R��o��]|���8M�_�i[� �dh���/�eE�[�O��G�J]|1oN3�ݤH�C�'��"~�=�-L�gw�]U�H���W`:N�l��\!�[~�q$�� ��&�JW��Q������hB���R?����/wN�����y/r��B@�ζ?��Qsv�{��8�&�w�e�>e'�Bq�H���A���a�7~��:���ݾ\0�?*,���W�Ԙ0_D#��}i�O
>�t�������!3S(��<E�v.���AD�f�*$	� Q������(��(<���|^"]촡���V���-�1�#��=9�Թ��U)�|����gdd=�HE;��|�d.ˍ�|*����v&j�2xJ�A�^�4��SV&��(ѯ�9�]*n�F,�D��!U�ߠF+��-�d��3>N�|>��n~��������R5P�C��ӮI�t� �萒1�g\E�,�K⁅�}%������-���xy��G�Ҙ̞��2}@Ѐ�%k١�"�;���
�>ta�	����L(�E^����$��ᗉ�\�����;�ͽ���e|��Ԧ��;C����t]�k�������0����\k"�f����[G�GlEnl�nڡk��.���>��h��83^z ����י����\,9Ǧ�N�q��B�Xj���>f]+���!���Tة�e�Q JW@џFj�ƫ������!3��v۵/���pՅC��\n_��867��"��L����8g��]Ce\�'��{�C�:�@��N=�B�Jڅ]� ����;�`��cl�a[]��0TO����2mh>"ZܗYKQ��X��H�U��XqK�~R��EF��j���2����hr}�궥���?�̒5�t���@p�U嬘-{�~v�.
F�q'��g[��~�:�r�����,֧&A�m�M��L��ā&)Є����HNo*?��&����
JKE���x�
�@�Sպ̀ 0��?$�<b�k�Y����`�⚴|��K�.a���cU8�\�C.�74h��k$��Yi�{c�����ƅ������ݩ��.��	�z��\��Z<����llڣñ%:Q���/)����0/q*������IkF9ϗ׏��k�d�3rg�F�� ��Jo;��2����!�7�3��I�	���V��&}��X��_����R���C���ma�;��e���yX9BVp��י���7D�Џ���b��{t�bA����-*B2a,���n�t�W�l)y�qQM��<"����;�=Q@�A���	�Qb8�F�\,-AAB�U�_1|�x���.Z�
 "�^ЍWs'b�4}(������z6��.��#t���U�%#�-�xV�5T
���d'b�׸��tD��t�>,�M_�y �����^5�Ns��tR�L�w�Pn79(�"k7
�r��[ܖ��_IrJ��]\������*Ç�Ѱ��(�ޔq��:HK����ܹл7�{��������z�{d��(C1���MJ̆�L�`]@�������o�֯��1@���IPլ�;�㞩���k~��,3V������%1��\�vpqBeO��AL�&�3fی[J����_��º����8���_��۴dpX�ڭ�}<�5�8*�ۀ���N����g���B�U>�2z����p�C�rÌqW��W� M�6��iB���m���K�2��|�x�]�����SR^�T�xX\IJ�rg9�M����1�R۾@\~v{� $cV�V?�U�%���R�^{�N����\�L�C�ϥ<���1s��e���[��S���V�f#F�����0�]T��/}R7�4��Vp`���n
e]����A�v�ts�#����(���j��d��)�2����X'd;���,Ca��dP��h���T�� �]�)̏��o2�4:��]��m���ѱ�	`���$�zG����!еs��1M�i�􆠋��ڳ.>rj���c�y�3s��55�L��J�ʁN�@��Zb���4��}J�yV��眧:�:\�fRݣ��3��"��0��C.F�J�O��sL?*�v�M\�݌Ʈ�B�ޘ�����ޓ%R
��J�&��tS��?2���`#�*�-_�LV����������:�T��Z��lֻ��8�G��'�=�5��
ǣ�[�\�Yuμd��\rO�䉝��(󫌧䃘���jZ�c�a���}��&i���k{5��̨S�ܭ�u�y�����¢?iH����������j�'L��F�#�~�kc6�K}������L� 5��o�Տ�������X�����a���dQ��Mbx0���A�!Đ��kSw�����<�EBJPea��_���<Us|1A��DǪ�p�����d��8�U��P�[�Wz�}~���r��OXѥ�0�y�f�����:$4���Wa$�W;����QV}]�V5�i����B8��Cڻl'���@
_T�^O��[ޛ��8��QO�� $��r��i�7���gZ��n��G5�~L_Z�s�*��
$S��a� ���#]�L9� G���Pi��f��,��ysD�;��1K�aF�W��Z�Q�E����<���Ɛ��V���C�!+��v?��\��lF��C��a�˶�,�`�c=�6
�@�_6SQ��H��$:˱��%�v���m1^+b�BpN~��>zrq~��/��k���-�>#?�f��jq��_M��4��f�M��8�
�L\lF���ɮzQ薑`�Ak��&�����h睭BL��1h"��:�X�t��2���l�"O! m�Mn�qs��C;��D�;I_%��_���)o������h�Z��c�Y�k5>��f+�A�ih��k��� ���_rr&���MB��J|��ư�Yõj�
�{b�,���p�K����G�j�Y��Ӱ��~�]N���ꘛ������쎐��%�>�����fꬱ3vxA&��u#�mz��y}�-�<Jl��]��*.m���-4B����'�6�R�uZ'��l3��,α�n<��j���,Cz]��(���8��_n���5�wT��'t�c	dd��pR�C���]d�LU�F�
�J@�� RC�[��^�6��.�%uJ3�rs���l7�BGï���z>tͬ��[_"��|�T.�,� R�`�I��fL߻�f��N�F���aEC�co��n~u/�t���vO8N�o(�H�Z|�*�qG@'G9m�`7�l���	w����/ێ[�̡y!�grU�7��"�(?�&�?��V�n�:4���.�yd���_�  �4��C*|�|UPbh�Od(�7�w؋V���U:��}�>+U
���Q�;dC�HI�R~hD�U-�-�R�v���D��'�>����_�ܭ���H�L+N��I���%~��ڮnc9�v2�I����2y$��E�1s5i��#״�\�GX�E��.*T+���IW�}�߯P�Eoc����Q�^(���'��p5�Ί�'��G+@�dq`��v�J��O ����N^囬N��%��܊(��YH���Y�Sͱ(o;��y�^g��Q��~��S�a]u���Ss����5!������ǁ����8���`�㛄1��X���2�X|�7&:�s}�iۓcs�G�����Wpd��.e�\c����h����m}��!@l����wԸz��گu�\��:��҇Y�/�7Ez� @����+Ö����p5N�
��aܱx�B��wqS�U�S�%Q���R��K�u��U�bC����e�b������"zyQu��G����
��;�����W\;�����^IH�oq˞N����i5�n
��+�= �>aD�u������tʝA4�������_������ê��E��j���y�f�{��b�2��M`�rH�Ƨ�u���oc%J`����!
,G:"�x���
���]�}��T]�Yh�?2}�q�U_�F��$�W��vx��$~?�	5��L��֝؈�b���vE�K��^/�KIL��g5�*���]�Q�q�g�.��|�ꭧi9Թ�H3u�Vk�T�I��UkՕ�ⳏ��
��ڃ�9�d��KS�M�R�}�ͧ9D�<�ߺ�0g�b�Eȅ���vZ��\��k�H�;���j����W����7�F��==
E��v Pi��K�b�8���Hr�V�P~���������i�"��A�s�]8��gQ`Y����Q��H�H�&V�&�4�Cd;��䋽/Ө���5̎4lj-���o����y��4X9����Ug��$�Є}��F8,��>�]�k��H�d/2&�||*����鐝M�i�d���˞<���ɝ�b��9:��N=��v�&��A��n}!Q��&�f��m�������,���ac���u�<Ƨ�P�g�g�O�]�8�����H���.<4?Nt��H�srFp����DJ�y��\�j��b��}L�Kq���! ����C��TxjW���3p7i&sb�k��JM���wtf�E���k��Ú/� ��!�2���|�gL��\�0EX3]aKc��dm&⃺}J���}��Ұ$��U��l��0�Z�ީ52���~�O>�o��S�{x� �N��N���'\�0�!D'�3�l��rOv�x��a]�Bdwb-�*6gG]K��c���ƈ&��݂	 ���4٩0Dv*�il��?�\j������T!:Բ+�M5�G-�X���Gm�
Í�?p�8�T�B���¨�c�g���-7@(	�:c��p��.N�׆��`���a�=��K� &;��ž>Z-���KG2m!���n	��m;�/�*U����޿-J�{;ld<p����pv�U��ot5��Ϻy�"7;��űB9�*E�kU�y�,�B�=i;*I`�p߯���93f��3A!e� �t������8�F�fyNzYߍz`
 '�SU����S+�K^�RYf�z"9c����T3��U�D������<$��>"��c8��R�@��b%��q�pH�!��ɵ�Թ�0X[Ź�q>~6~բŀ+X%'�=��>~=Z	��V�*��X�q.["y�v՚Ƃ
��4�1�|�x����t2|�ʶ�k����=/Wz5�c8�mk8%o���p�U�_P�w�H0U,.2�7��^_��kI�\J�(M}Vj�S��Me�3����3!���G������4�#X��|�ـN�&п�V:]
p���̮E5»�c
���6x^��C~�X�5X9�	��'���fcFX%��Ѩ�&���Ɉh=�{0��n����H\e��kqSv�6��{>-�C�Kr�V5�I���D��N�(S�)�l~%)��#���2��SW����=�qJ7���R��}��縞M��W ��1���>�Za��C˷��~a��~�í���Z�g��,!kH�$���0�}idn�*@  ��F�B+�w�]b���)��Y�����ٵ4��c,���NB�����F�G����4*H5�F�3��ɥ��u����Qal
�}B����{ [Rϱ=1v�Q��<�8r�ޙĳ�����ۺu$j���}K�0��C��CbV�4��s"�2+8"�	l��^���}�[��*v�me�P����#�h'F#��<w�wa�of�1�T�Ex$|; .��������̃�%��9-{V@)�u{�Û���
BҤE�`�i��G�b�̂_��^�~*���½)�_��������ְ�hb�o��U^�IxP[	��8Q)�����`8�r�^��q`�%�K��Ԕ9�)
ov~���cB��	-�4�-�2�S6�m4k�'&�+�RHa�l~��P�6S�bҘtfL�������E|{ڥ˥�g���W�f��ג���c��Ie̾�
`�t|�����lX%͎��_,��#U�^-=��1�P��������Ԃj�/8+IK���9�����9�\b3�0Q�=�ݜ��$0�1I>�i��W� �t�MW�d�wr�\�2 �od�t�K��*�VZ+ebV���^��B���<���>�e�0'�B�ї[�������h����:`H+����cĔ=y},�(�'׳������Zi!�`�	v0�Bt�*@��#~3��Jk�[���Qc�6�}�P��%�(�����o���5��_@8|y����a���.�=��vKˎ��ogI�֠1L�LIfK�����.��� �NQy��?��-��Y�æ�x�{@�(�W-�+Կ�$��՟ 2���~ґ�u��j�坁��|���i�K�v��d��;`c� �d�`߬�3=U����t�՛@��h�mHD�0͛�m`g�0��[*P�aBP�iyJ���˦z�70* ���A��u����\��YZ�vo��\�Q��ĝ���|Uޚq�0 o��{���i�W�-�B�^���Ĉ�����0Ӻt.y�Vr�ɉM��\q����{����1�xN����̎'D�
���HpN�n7P�ս�i>�Uf
���#�
z] p����(4'��J�W�R�.�ׇ���Ko*jxP9&���	{h�a��_M-Ƅ����zV�|��~�����҆CA|�lM��e<ݲq��.-��M�_ΊMD�:�h��_��(-�Vp��KVk�N'X;&�D�5��ʖ����qtVgYA�Z�u@�||�cb&�z�4�!��i�LQs�9�������2{�,B^2`P�&��&��Kx����`b~k����k<c�{t��u���ۃ#7�<멅�}o@=�ɧ�����F��T��K� �Jt,���4�hJ�.%�O	oY�if�������_����jF�qgh+(?���%�W�i7F�fj�n��|�h���� ��2M�h�WCRE��殅!�	?[w���3�"�n���i"k��l�&�̯R�Z��昖�Qf7��xeB��t�w��ͩ����΁���h�!����.g����ՆX�m�%&��A�F���/�P�/3w��Sڈ
��?�y��21��vh���Ew����4�'U���Oӈ�Ȫs=,.�
���ɛ����U
��S���*7L�����1��{>�KM�kޭ��v��̏0a����f��@Ĩٯe�H�a2�Vs�H&�ca�a�f�����}3@��D6׻�=�g5�i�.��O9룃���"?):��
��tW%0A)!���� ��(����G~^�9]�iu��T��+V^	r5��`�U �����f=���y-4�Q�uo`U8Y,oѾ;OBrT�}:.=s�ү?\���;t�݌!�Čȏ/��� �+�}��:v8'nY��g���=�t}�OI��Ԭ�?^�����=c�'�'�7K�ߎ�Dj.s��:@�WW��ã��ȏ���:Th\u<�V&�4�D4}k�"�p���j��(�a[� #��4_�2�Wƴ�K"+�R��2hz�=6��f�o��r\�����}P�1�v����ܞ����8M5`����Sڐ��+?K�C��ׇcT2ϧ��X�f:�Y�ZQ06)��Q�	)�y�a�!��^�\J�-���܎y�h���SU�5��T)-��W��hm1YªLJ����Rԓ���$p?k�7��A�V���$4�¡�,�8,�Ҭ�K�8�.�:x�� �2ݣ*Vc�Q�c�w�"��?���#�9$s�k�Oǔ���9�_pl��y���E�]z1��/�a֨U�$R\9�����O�?UG�����+I�
=$x�/�o��ɳ�>/�=+�����)ԓ5iB M/�b����4]#ް��w~`�Ns�;w�����S��8��Ib5jwEj{�l��ir�:��=��9�&j��ߩM������q��)��(�MG����u5�lh�r5(ahܬ��*��jN�����y�&�������e,�=(`_K0�}�B`��E�H�gr��ω�'��c]K��W�a�����ɨp�g7�A������9�F��Bl�-��k��g�ƕ�8��>�4��Q�S�F� 
p��E�<�����_���PE�NN�y��)���zP@өu�È0�͚z� w�Y�j/h\\���t����x��׭����ox�G�ޣ-(�Y����3F��;�(������z@`����ԧ;Gsf>�cc��&���%_2��4"'�^e�}!��$���^�2�� �\e\� �D�9z\I>i�9�a�����aa���O����łU��E's�_��C��1�Voxk;Øلс��ܓn���zR����-	���$���=!���O��N���ö��<�bۻ8�:�*������we��k�]��
�p1�F ��?I�0�q�N�^E��ڧ���'�/
�lk�Z�Đ�Ek:�:�_��OYbr�M�]�M4 U�x��/6�Y����YKA,I�e2Z/JE�l�d���"!� {g���m���C-`oS��(�����}r�B�s�Y�ȞN/���h��^A5����6�죚���L��2b��ͻ����]�>��|`�!�}9�y*N�ģ�\li�'��%ZE6
|^W�@��a
�?��e��`U��K�~L$E{bI����b2�/P�������={߅���t���i]�l���*zi*ny��D�Ծ��6��-8��;X�j�A"F'�-@�b�B6PԄ�4Q3�Н���`�Ë����G"����)�m�
��OδB�t��\�A��M@��Б���o�f���7.���?7��\��K�O*�����������4��gYW����O�^Ii�!�>T��ʎM�o�Y���YE<�H�E:+�'��M�G�-��}��D�;�Y L�鄅xsL-���	�#g�	�on��y��ڐЮ������5��R6���b�VP�+L��{��k��r6er1��ܛ�Ss�M�JƹT!���r��}��9�!���a��#QOu-X5�Y@B֙��n�RS���Aᆚ__�^j�U���j\y��ރ~�f�fͤmb��:�ٔjX를����Sl�8�� X��Z�o���lp��Z��2Ѩ`�aĮ��_�j���
��0w锴q&d�,%"Yõ�(��^�ɝ�(�ܦ�
��NEж����?p	SpT밢C�)�9.5�<'��ǮQԑy��Y��m����O���N��1l@��	�4�(�e�� �!{K�hՆ*�
�sBҧ���`�>��/��ʐ5h9��l�ˎ���E�z��Y�G�9�	��`O��?����8�ΙswK 9)���{7��UaJ�e�ϐw�W�\>�2xp�
�!X���}�����	w��c����S ݛ��dY+~䋼s���n�c�3���J�w��n��x�oh]�;��J�PC�R�
f&��am<J�a�W��)Wc��E�t�^	!^s�t����+�����.�Z� Ca�Ei�)ʧ"������ ��v߼-��X��a?M���l�{�o�_b�`C�^[�5���סni$�q��/D�HجH��B��ʠ�i��T��a���+.5a�2c�89�7��h�*h�(�d��C�Q ���'�KM�N����@�B�I�"h<�M�B��!�y�W�ᣧ�7�0�o<��r�t��UN!;#c(�5�4��?߉��5�q�n�罆�
��}\��4�JCp�ӄ�Ͱ��V%x�Q7�/�S O�?R�׹,g��O������+&�&\|�c��΅�i2��(����r|�R5Oi:�']D�$��Hc�ȩ�Q9�������utu���>U*�\���f�G��,g,q����
���[�;�sS�H��W {��R��+�Kf�s������$1���(�U�&�	:K�����]
�l�͠�6�!�7,��s�(5̅�7�UU�<���sF�TӨR�a 2{�.;�M����51���M#����8���&��1_�y�C�5��!����-u	j�w�E �/����Y�|N�s�j~�ak"�|�4ه����d��|�w!l*���t7��ۨ�������DH����wD5�[p�B�;+ѩ��
�~<��:㭄��~���\� �c��zj�"�[���k�~F!�֠FKl)���{�������#
���P �W&���#��ăQXf(IMmO���s�f@����1_����[θ�v"��>�<[���D�n��Q�Y[�s:s�)��=vښ:�J��W����.a�A�-9j�uw)��߉{v��;ç�u��r�q�"�����JҟdzY!�`����C:����ҙ�]��Gc�e7-X�d��%�yc�dHΗ'2��H��!��r�i2.',��� ���ո�v�o���$�v	K��<b�N�Z�,&�8ءS;E%�isڠ�Y�7�A-椩���7��W2sp�yO�fܪ4Χ���	�����'��O�I�W���|�c��s}-�x�?ul� z�K��n~�M0�mߥ��R��;Z��4��[I��K�0U5q�}ӷ�%�W���p�%�b���;7��G���cD8�p���%�)�9wȯ����nyޒf�t�%����4��ϲ0C7"�#��ܹ}z����s��x�q��g�ܼ4�}�a�`�_��X9)���l��zV����D���q�8������������6c7r��8Yw1����+���S��{>x�k��9Qb��[�����(֪@L�]�k����d�f�|s���|�9�-9���.�7O�Sz�f9Ns��3����	����?�� ꍜ����%�@u�`���N�|+�Tޥ���|�~��tQ���~^5��c��/�k��T�|y��)�m{�B֑�h���(��i�]�5l f����{�c�
�*E�D��ui��1\�Zj��lqm
!*��\G�� �E@⡝����:����d��	I��������z �Z2k��9l�DM,�t��tRihE�u}D�%�2��7��F�p9�\���u�G��q����U
ir�l��6ϗr\�.���mm{��X&[p��������j��P�w?�-~����H�) [4�$9�PS$�8@O� ~��������%�+�.L�Uy�`0`3�����b��`����$�*Z?sV�r�@)w�3�*9�����(�ٺ��HA�ѷZ����n�Zd[2�#����P��ȗ��i][��lo����{��4��R���߽�����R���t
��c|#��
㌼8'՚�3��Jsg�=��:�k�Ļa�^�m��J��C3?.l���
������n�K��m��4��Y0NO��Mߦ�ɂ"��(s�_b�F�`�!�ym�,=ݯ��;pHMBd2.8���lV��W��c �9�.ϫ��sOO��<��B��PU�}g�� t�ϱxvk:mYd�D�4$�I����d*�d�0�4".2霂��}��p�}�"��X
.QqjhE\3�v�K�Ek����:��|]��Y\P�rL�����%�����V��E	&�8�Lo� z����#�'�;:^`��bF�Ni���ј��z,�W=Bl�{��\�w�N<��`�'%o��}.��w���j��~Lr�!Xu|sӭ���b�D���p �ƃ�;7�y�CK[��c�±tX�w}��`L����Kږ�W{������h\�XzL�R�����r}IK���1
W2��χ�nD�qZ0��,��m�c����#]���������k'�"4�k��7 l��H�ź���@}^L��D2)�����շ��P��o�6�7���#��v��]�-G�@�Op��4]�	���.�9X����<����t�r����~>c�9m�]� "��^w��;���,���v�*��q�p�1a��f�9�Yep� F������h(Qb1?�Wb���4<�.��1��b�V�@��� �x�g��eՌ|�!���Kuz
��������$���"���f����#�効q�w"o���b$� �f�=��LZ�\'E�8e���gR��UB�/�fX��34�m�sS�	rF��@��q</@�3ԁ$������J��i��L��$�\�i��_o�Js��	+y!9�uK�*|͜�P� �&��#6�ߦ��U%�D���a��v6R���P�i�L�^p�ת����ߙ\�g��J ��n�7�t06��9e�5.F���'FRi;c�����l�^w���@��|J
rj��Aٝc���Rcb(ul
#��(v�×�	,|Y�f�rd����,����w�(���%��Չ�פf��|ԫP��l�#oO7Y�4��5���y>y��[^�o���k�iC�^�~tdQ��
������ߜ��yn��}���$_T�4�֠|TW�0
f�+'�W7E�hI��\]��[wdݏ�tMT�kv}��!t����+�8M��9i�c�	�N�&"�*��|xhz��aO<��J�'5��	_F���C�w%���@rA���0�f׆���QR�,tW������xj�vW�D���w�du� 4����0��ٙ���oq���j*���?�)G�6���\	:x�숺3@��,s=�z
:Ԥ���7�LN�>��8�2\}����J�坸zڝmp�
��u���2q	���1�U"l�t��ϛ���2�ťچaV�P50�3㖷1}�J��!�wuO���J�-M[�ֺ�x��+�Y�Ͱ��J��	�mK�B^�"���
�
>.�0K�����J$ t�ݤף�+o kXU�k�0���eF/!S��g�*��y靈�(�+���o�G���(d�çQ�S��`+ WJȭ&&Ӯ���	�L�h������k-{���<�w^ܾ��8��6�$��K�'���[��l���*yl���W��;�{zy���ݡ�V���W�P���H��4������[@f���ǆZ��g��7h_,�ɗ귍�Q��Ɣ�h�/�D���{��\������6G�����2�#��g�^�Csk�"
<��N���AK�Z�k�HWX�ر�ǉ:�~�h_�K��U�GB�x�(`����%�l_�w@A���LA�gm9�i_���0���T��˞�"]r�P�i����X�VRK�+H�Ϟ�_O��W�P�&�P�̙����߰�9�y�u����<�Y^#0t��N���%�օm%Z���~�G��.}�It*>�T?z�� ��RI��wٮ�u2�J I����H��Lw�]|�.{�۾5^5&�Mn1o^��H�8;��=z���p�u;��O�*�N��a�y
[l���{���_h���Ǹ#|�S|�K�o���f���ƅ�
)�%�b�7����l�\���r��Jf~.@�JKCmI;-g
�rŘ+��w�n�Mhe6����v���MW�����p]졊�d�<�}6i�u�ꋿ��@id�ʚ��� 
f[P�ڣf+��&Pzx�����q&�!Q٘���y��[硛�ͺ2�6���B�� Ps�w�Ijf!9J��^�;?Xy�)ڷ�v�}YT�!��ҧ������������RP{4��h-���2�5��=�A�����d}f ����uMQ�4ֶxo�}P�Ⱦ���E�@}>��� ��ĩ_�5Yٟ��`�S�U]G��I~�aL��:�{�ۧ\޹���L�RnQ'��|C#�������%��\�=Y[C���o�3�A2�sdV{y�����/UU;$x��8��;=:�<�6�k*�-P-��%�3}��͏<��>�����\eX�Hb�����3��;�K��|��	s�>y,F�k�t�(\?`%����u�?��*=U��b��,a�HM�U����5�c�*��<���b@��ճڎ�Sڽ=c v��)�Q���l�5��>���8����UT�U���5�m�jQ�J����\/6�5wFq��{�S�R��E:�V@h��Gd��!�e�!�Z뒿�Sּ�\^�����E�H\�x�{���!�>w:��F�l>}	o�V�	��T����_֋%I��1��E�/�<�8�`������Ќ�K{�<���2��IxF���`ʊ�e���U�-X�C��6l�Qw7��J�P�a�2��v�8��"<�zs�w#�2j�c���sY��$[X���R��\�m|�p�}�M��dJvv�L��솗v��{���p8��#����y�z�.XT�ͳ�
C"�n�7㓶Q��pY��%�g>M���}@�	�'��fž^#�R��	�G7}i0�e&2,�9�J�pЋ!���E49D)�Q`7zɯ��j�[�gl���LS��;%��������re�1�6G�	��#�'9"z�xy�If��5� ����-�
g���i��Z�S�y��~��dY���c"�����1Ջ��yF;ҳ�2N�4Hgʗ
t��T:�E�&�����F x2�$ ʌ���g������EY�ݯi�h�^�Q��&[3P�P%�*x�m��K�l�ˠ"��q
0�r��楴ٰ�D�hGT�SC�O~�������4
�<^\i�`V 5}�L�%�60s����&?p|�N%��#I�\'�_r�GRwN}i�
�Ui��?�M���Q���*�(V����T#���O×�G�>���;N��i5�#�8�NJ8^��?�Ouun����|���@a�����$PemS��B����)�?�9t�ޅ�g�}�9��?0�N��а�>���-R��Z�G�'Xsײ��>M�[�tM����2mF�U�"?���a<����j#0}�H$^?nr�Y@Z];i^p�*х���؝����B�ޞ2֟�n�+�${��3N����WH��dK��4�ou������f����j%\�
팵���"r�խSV�a�3�ۙ�x��k�&�w$���C�^�V~All
���Z(�we�ĵrh���7~%?��5ѐ#[�HLώ��xmү<���[a�f�EK<���_�' ���;�<;�N��omZ*@���`��m�>8�g�'A�
�;�����J'�|1�}6��4a�4�^�p�V�Fb�� u����:���R�+��~����A�ʕ�l4Gې-~NH�v)Q���V)
�G����5?��+
��5o������ʁ�a�~�~��-i�=G3��	�G `@ء�[ �j�
�Pj�j]�Cpgޥ���o��`����ѽ]Q�w折�D�X�®G�����sF0��u&�e	W�	}�Lл}�a2���j8bS����D��J؛�w"�K�V��f���Z-��Tg�Ó��dY�.8M(�ѻ���ڼe��?�{��d��'���

~��7��·q�a���j��L�k>��8��s��ȱ�
���t1���~>���R��?5}�N�F�5|l���eGnP���b��)���r����?3�<�]���M.�? 1tD��(��h�U$�H�o�N�29�M�]�}b\��Db:��u�.���R�;"��n\5�� /쮫��u���g�����	�lt�K��]q��q}�|,WZnˇp��� ��n_m�2z�(��ȴ���'� �9�!����3�e�$'V�+�B�����z�`h�|�?�
�TzP!"�界��Nֿ�Dg��ԮW��_T5��p-ܝ����������c���.��`���A��C���[��ٕ���lz�*�srѽ�IwF�~�[y	E��W�'Bk�y���D4��q�p_�C ��k�	bjJ�h�Ά�ߘ	1G��H�K�Ѹ0]�Y8����מ��,�[N�rS���9�}׀�[���ny�f�hL��_���Wg���V!f�
g�s݆
t,�������n���=�"��'�R!���N�%J�å�M)�⎕?�;º7���|���U��=�(�	G���|�^��SY��ˎa�A��mEQB���]�y9�m�	˪0:E��%���V���0���0���T`��:�{�$�Xt�g�~����w	޹X�B8u�����B�Ju�}����M8��'�eC�ū}�<?i�&A��d��e�d��=u�I�����*I�/�uЮ���La�-K��;�^��8F��Y-�G&����-]�s,3l�����)����y웦t�4,5�(��ׄM#T�Ԙ�m���p��������!�A�5�iB�*"���{�U���pq|CԵ�
Z���շ��	����>f �� �j8}��x��?w�l ��<`F~����#E���,z��jR=���}0M&|�Nqjɻ����7�·���iʄ'��0�\ZF�ն5�f	�����rb�6��t:oϦ�%�Px��1��v)�n{%���c��h�p]�q���,s	������k�'xX;�R�vG�ocl�@M�y����] $6�랉����%in R��}q���Z� *4�p�5�0&%�,���n�=0��azY�&^���%��=���/Za�:�1��.�àL`�~�y��w��)��HȰ����
��W�F|-�1�@k:�߬�ț����S����v�`�(��J���\���g� lF?J�b{��S�����B32�=���p�V��v���}�!�4tf�8��]>�v]v*Y�ޚ�6<UN!\!�'*�2_��L.|i���U���_�&T��O1��L��������� ��)Ӝrf�reh"2gi�}�(dʭ����ەq
sO�X�8�PF�O%R���������LфF�[�!�T����5��E�a��Fn���imO�0��L�E��<��萳��B��+P���ǲq#�ؒ�Qĝ&��r;ĭ;y\�U^���/Tf���l�^��A�q�=��\�dc�7o�/4��:/$��dZ�s��6Ir��r$���%��aZ����\�"�:�m�)�l��<6-�>���_e荧�}ႫB��bEx��v��I�Ǚ�˔W��#Q�5��6}�%�����pl��|����<e:��F.��dN�Y,]�K�BDg�p�˪��5�,�Z�=f�� 0����L�	�4�&��'G�.fE��|�knt�j���RH
�Hr�f��R:X�n;�s�
�&y)D� }?������𲸧��ة�q���{�IS��|nr�]�+�xGy �����[H�I��I��0��В���S������=E���kQoN�Vƛ_�Č�7�x[*[��H/yB�:��^��5g��s����;�9�Ϭ���[q�s�G9[��O��X�dm?Ҹ�0�s�E#��i�wE4�Ə:����G~�F�lh|b��T�.���Q8�}�0�O*M*�z�X ��r~@�����9��2�"�S%-߉d0�E�޹�����3�[��jυD��dƽ��d��p��]p-&N^\�#�R�+3�$�_�������|�V� ���n��s4�J's�����A��[K���X'?F���R<����P@Fh�dyu�I%�zc�H��J�a�U:���\��K0�o�gWf��XR��-�y�����&�m���4g���L�ߎv�O'��,��V������6���v2Ò�*�ޝ�@����7�Z��k.�\�I��ZK�wH�>-��7�l:�1"Aj�ے�C.5����?�yGG�J �?�s�n�Qxp�s7����q�,m�wi;�}r��h�Yu"U�#��;!B�]#>��ܿw��H��(m���g�Ͱ3P�;�� ���Y�᳷����܈/r��,��}K�:i`4vVo���a�(��>��9ڎX_6�T����s6�v'W�:mH�����AOU�C�C(*)@v�fV'y�ꗎ�4������BLv�پE�`���8�5��%��{ݪ�;5�N<��t���x�V�=�LK�r�a��F���9:�f�">K`�S�k�J�O�`Ll���ٷ�otG��u�y���g%,��oa�<Ɩ��-�QUJRdZ"��5���5���^b�P�ǣ ;]ͬ�7ш�I�:!�8�
�ⵞ�*��Eu�S��#��=�~��ٍ��Y��C:pBҌB��g�i��u�%ח`�X��4\+@u�ޠ ���[p+����m	z�e�<��x�G�U�Z�|IX�;s�6w���S�.�#�*�i��#9����rN�}�ݼ��y����]k&����+1�(mL��D\n[��!�Y��(w&m��1���}>�Q��)�>�͔o��M|�1Q��3�o���|��A�iVj$���V"< MՒh ����M}��Z!�O�C%
(�N�x]Qj2�i�}�ox�N	�dz���[�B��!�]�Oe���i������ia�i��t��Q ��8�v�+�iv������>�����9&#�F$x"���	�5I��է�u=3�ab�@:��7W�p�x�@�Vڧ���˫�j����/�˔��e�zN����I�8ݍ֥��	՛�2oQi�
RKϒ�,`��Ę]��\�H*��0r���p���������ܓG��\��PƼ��j/�._�d|���:o��c>QZ���l9]=���p=G�!��J�^�m\��%������� ����HY��?�V�r-mOt�Z�AQ�=ci���ПE����y'�Z4��Diq�J���l�j+5	V�I9m&��eF�D�j��a�OK�@Q��1�^��R1���{�D(��w)g�)\u��6Y��^����S+�bJ���b��9�YNB��6sK����'F�aU2cRp���N=�kY�Z@�V�$��:��9-J^e���:�/�Գ-��{��Ǔ��힥��c5	�pý��w��G��ퟅ������*g���z^ <)G���rT��w`1r���z6bY'"��Ĉíᠯ�-.p�*p�:;r�lx)��7xW ��Cc�Mj����5(j�!u�b�ʖ���0��}�"�gi�D��h����8{�E)	�O���AZ�� o��A��h-���sU���ь�M(�a��V?����o+�'?�xLՅ�*��|IɌ�3�*z,���2������馿��_LU����/�4�8&��8���s�<���{e����� �2�Q��O�i�X*�[X�(RO?Cm��	m��
2�ƿ`�G��S�#� ��-��*&��h��l
l�@�A4z�vؤ1�g3O��8	�]��_Z��>�5�ږ��"���'���rhI-�܇����<ʔ�a�N�?���O/��sȚOI,��U����*�" ��[x��D��t�M�j��ˀC����9����>W�?>I��=��Hމm�g?�7���vqK�A
v�	M����C�
u�_��c�S&��m�á�tun��iFs��*c+b��爑	��h4������=\��}D�^��TV0�����0i�"���7f��Pm�%m!ɺ��WK���u�B	UdK�ZU۾Hh��$��z�WD����
��8&w�K��tr�`x~�M�~D�����b�A��#xy�ZK����~7��V��P����*�?���_�:,�D�� ����?2��07�'y����^F����R�ӽ=��R
��d�5���Ş���(
͌ł� A��8n�E��Upq��ݺ2zů�tZ	�5u�e0v��P�/�#;S���_���ז-��b��G-4��b1v_�d�3L�j��',�{�	����F��U/�'�0w~����at�?`)%4�R?$~�b8��gӴ��>�o# ���c�|IA�F��G�����>Эr�nDfa�Qp��;_�i��D��#L��@gG�e����)�����i}�2���&���d�MԗC�;�8tĞ}@��%�s%=y�E��0�8أ t�#U�7Q��yc�i����Q��knJ�7�������ծ�0Pfr��3��"o�N�r�Q���%��nq�Z�2�k��&&sh����.��+�`Ď��J�����\u}�ڮ3,�Y�;�!���"M�����[�^�'&yd'��#/�hoLp�ub�?�����}�[�2�����.@7f�n�Ŕ��}�O��w� ol�p��"��C:��&�B1N� �'$���~CI����5z��M��8Ү'W�O�=��ݵ�9��!�FSj�ԈU��\�z՗�o%!���$�	�6��]̶5�K����3�j-X�{���
b��o�s7���o�V0r��ݔႫ�[�8�9�@��9���Λ9�H튒XM|7S���_&��hΟ���E���Tf;h��d`'Ƥ���&�}X��h�ȋ� 
���F��{'�T�2Ev8ۃ�bŖu�-	���b6�0�k=&�f��&.�S612q��%�f��\�cz���{r��h����0�n#����A�)(����b:��?}�%MWz�zs�z������"(5���=������|( W�틿2�B��p���}�߷����flF�y/\z�!��neY��u�g� A=۰�Ksk����K��ؙ7O�����YG+����8�T)M�c0�S'���IEK���Ŵ�w�j�ـx�����x�L�b6�1��A<�7���ͦ����\��E��KnZ`�� 6�K�~6�H�����z?�Nn�!]��a�E��?]h���v�������Y��� �w�&g�V��������:0i�E�\l*k��}�����[��h�zG��0�e?�RGAG���ZWQ?s'x�gOI�ᖐXE�H���b��eA�)B������T�3�����S�v�� ��� ��KQ�M �L�8k�Soq��jh[�&,J�_w�c��ɓ:�6Dɺgs��&���e�����)�pRA	����hw+�Q��:<O�s*���#�}�y�z��f}B�`���[-��B���Y��$P�Q��D��8QrU���;(M�M�iE��d�dC{�<U�����&�RzS�"��9�,Fv��(��D~RWڂ	ht����"$�qu[��u�`{b�����X��	���mE�u����(7��3�� iS�[��4�e����˺�O0�H]��ч�a�w�3�UZ���w0wX
��(��7�2�r�0Ϸk��>���^_"��<���ٶ��2��l^�n�K ��?;�p*�������\�e���*6����R꥘�I]ώ�O���Y��~%������C��by~�$����c��JC�pn&�o��/t�?��L��������/��迆��s-�~^�ޗ�b@ � vL=����������%�9E��G�A �묰d��{p������e~*t%]16�����3�s�$�S�  ��=�:s�1pIÆ��	|H��E�������,�����vWTUY����A��qn�V�|��pT����z�ՌFf�CVk�2ag�u,�A-0'd�"H!���<wZ_��t�8h�����5�`;l���?Ef��-1�n�w ����bFݎW7_���]����^F��dŁ���~�i�,����A�5�d��T���N|;�g�'k����K��t���@�����b��/����w�	o�̥����yr�������Vi>���w{�#)�^k��%<4>n}�k�҆�����3�Η<��������<�<�3�%�j�ݕO���"x@�K�H�s��G�+���
��-B���r�p8 +�N�~y s^q�!L��g�&<'�q����)��� ^�2h�cGn_���%5J<(-px�Nħ;q��$���>n��o�Ka������߫^��T���<���"C�Qc�}[a�	�Cf��|�����2A�e|uy�9��W��D?s���XC��;ڛSv�.�\?�TϏ� h�4������'�P���Ga��6�������4�i;�{�ܒRDH� ��GvJ�]`n��R��\9��_�fr~���Ff��Ϧ�ƟK�/N�5��6�gwA	{A᪞0�з4C
�q������U���{�K����\� �� �p�I�?!l'�!-#0q�:����G��6����!��f���J���װ���L����ߓۃ��_ƽ�Y�<��:p�6�\��|�)d�d�R�wy�˺\�ߠ�Y��b���A�!p�����)��?e���r:���޺�+�%R^T��	{AlRHQ��@�4�Xkr�ڰ� �y
��pc]�b��ȉ��:~�nS4�/r�z�S��@��T�^�XP���6��U?�L��u8
sb���[F�
!�C�<��iׄ�e�	Tqg$�-n�)l�T-f��~�[@�|����r�dB\&�L�;�M�~�n�X�L��.��]��V��:�N
�G�ձ<1���$�8-�Y����T�x����=AnHF/��pzYc�R9� 3���͈���V�E�����E$1G3wQ?�o��N�`S$��w�ʣ=|���<�Ϣ`C@�U��P�C�=�'����>�~�{3l�ƛ�cB6a��M8la�XL�֤��B��F|����W7&֞Z��:21�|I;fsA�)�Dy>��L�b�[����D�5��<(���8� ��T�ۉrL�+LᵳF�n��̮Rݘc:�<{��T�F����r�6�)��sؖ���<� �<I� ��́�Q����ǟ�����{�B?#��wT]��>�rE�^MeA�[��5��E��Y�?���%��,��5�U���qm�1G��ۡ���Rh���j�F_�I�u��c*LFA�Bh���܎�޿Mmu��%���n+=RVW���b�]�+R����K��W c9k�i�7�E���Gt&�C�{H�������������*hD��Ĥ�vWT(͌j8�#y5�cc!�mZ�,\�d�T��Mp3�F���*O��p>��QJ:�n�
���M},;(���i�f�k�q���ع�a����.�Z~þs�G�����	���	7���F]��fרjW�a�!� Yj��?�.�Q�:�a,�֚���,���Ƈ(>����!XaE�f�Rs�L��}@�"�P�������hh��硐��7d��N���]q�2��z���E�n�Ȑ��3��4j���:M�.Z���8B+�ƞ\r+m�d�Y'8?N��=M=)�_�w`�!��'.��P,��+�U|@��7h ᦹ+OW��w6�J�v�����u�Ff7*x�3b���|URÙ�!?|�@x�t���,�4���]D�f�������]�C������5�:�g;ㄣ���S�J��C�N/�7�͠��ǧL��?q���a-y�ZՈ�Bl��A��[U��S�|ҽp����~cY,��2�����.t���]��c�Dw5e���G(�@b��9��Sc�o���`x`؄4�Xy>9"n\�ȏ�Hdb7�]P�K1hN�z�Y/�@	�D�qe���ӕh.!�S	�@�[Ζ�ϻY|���u���'�;R�����-\��U�����_�0�P��A�4&���X:��Q��@����h��K�iQ��b��[�c=��{�~�s���[�	`��g����!fl�ǁߧ�v\�!�-�O)����.E����Q��M�.��R]U(��\5[��1�W��8��c�ΤA���$Q��W�ɹg@���&����,4��l��~��3�<y�A�%"8�7�����
y"8���kg���3k�}�,J,�ހ^9S[�s �p�z�������Զvm��7�ʧzG)r������'�n�b�PIkӑA볠�TB.�% �[ظs$XC�%���zߋ]�2�F^�/%���9_��ʹw���h�Έ��qsNW�)�P�`������/{����%��9a�q��L��7H��_����s�Y��y���ʺm����|!p�*��� �J�Fm���֑����DT@�z�^=8W�f�!s5j�72���O�)��?�o#ّ��Z�4��?ő�?�@���&��V��\�Mr�
��K�h�>��1�2������B�� 6�t'�ڸ�# ?^̌�RL�nN�ˍ5_�T�.�%�de��)9?��	#wpB���lE�
��Q�7de]���ɠ"Twu��u�t���v5�O����\�;4����p(dh<(�[5ջ�����fݏ�-�sҍ��,B.)�X�S��_Q�h&S�p'�/�7b�\���v�Du�Iz^���Tz��g$���.��_����x R�P������ֱ��ʈ�!�qa��4�Ҩ��}]�w(�.Q���նCD$Qr#uTH]����_4.[9�G��*�++�{�zn[���fB�reT�psam��i��c��ׯW��J�落��htf ڍ�q�h��iL�t��a@�[��eP���Ol2��>�:�)�)��\�B��Iѵ�h����I4</R�J��C�$
쩌'�t�̛6�S}���������镘���e�����@�����&kk�	�b���4��[���Q�K�IM����Q�3��W
�p�>�1C�y�ܶ��4���$Z�&o��^��3Km���2���D����He��]����f�J��(P��6t�I�Pk�K2�SQĵ�7}T��5h��X�X�G	�5��W:�� �[|;�4[�'A#fG�4W���>�t�I�&�9�,�KU%g}�jq�*4�\#-w��ܩƭZ�r�ק��~x�"�(At�.ju_2�/XC�n;��QF\&Irk�
� ��@����8�ɓL��gd4��W���4�;,FM/5��}�0�@��D���äL�@�<C�0#*"k6*hV�RV���w����pe�u9���ss��4�� �<uU	��7	�S\��%�x,���=k3@ã��=�~�N��uSQ�7����g=fZ�Ew��^�B��S~�ݑ�+8@&�V���۔��`�H��3�Y�^?�_�,Jĥ\w��� �	��x�4�Y^������!����-����B�P����$)o�{[�|�"�gzi}����K��t��L����,��&poN��Z��C����B��/�ޒ
��v���S@3B(( ���}�����R�2�$� �b�\aЙF�=�F��W����5���l�9��L{Q�W�㍠߂��}����i����z.QՀ�`~�-1��z�9|%~��a��wLזL�uX�꺼�[Ec�I(sꌂ^F����9�����<ϛ�M�8���L�Rĥ��K4 du�e׉��
;��DyN: � �kJv���j/��U/:�ӓ5U�P������3PS!��M�tr�?��fq֋:xh�-B43��( $���sx!�<t����R���WQ��:�'q�ݐO�Ͽ���P��ػA��.ͧQ��G�[���ā"O� FKO���'o�q�}L>fR>�����,��~��w�a؞<S�i(0�Rg�4\KD���߾Ȗ�-��ɖj�P�GK�큹u��NX)\3S�Y�+�.��%-\�WY��sSlo���^C�<�������p�\>;�\��4�8���?��w���睎/���QP[��P�^�'�׫�2Ҧ����uI/u5�n�5LG��~��|?����7B�+�RH�T W�UH���
��d(���|���&���a���0��缎���b2dQܴ��2sP�\��P\Pg6nlx�^���ઞ��͚�Y�.]9IM!����j�jb�`�㾧�ݵ�9�g�'�(�aHY�A�]�j���f6R������l��t ��W>���A/���^C���*�Qa2�6����3` y�9��S|]AD!�����u�5�ץ� X�\��W��G��6z4��#��� ��1�"��.�:8q[}!�!�Aj�ԠdK�����^��{�����1ct�!Ft}]�\�!��H�8)`�P�yZݾ\�ͦB#��m�)mz��it!�{�yq����X�\��rO�LJ��	�wQ<��;���6Y��%��/��M�4^P�D�*}lr�س���>�j%�>zC�3��\� �ږ������D��Z���Eǰ	_e��K�#N�e[_��}mqC�F�P#�J�e=�8��M����
C���m�%S�2h��]n�j���K��^�sU����?�9݈3�٨��\iYW`~��M���E�x���灵T���I�:8�M�V�4h�����e�e�C�z�ԃ@)k�c�>�_��Y���m�ۂ%��֬���b��OuxѭKot�њ�Y̲4z%�HjV��0n�Z]:��\A1���Q�x�Y?�lG|����6�!�y�>����
��C�1�|���IB��4�T:Kh���Ɉ�ۯ�hQ��b��a�_�Իw	|������`�֍@�tA�|�2�H�IؙKx+��ԭ���,n�9��|ݳ����� �����R������nOSk����
�VH�[)E����Q���:vt��`k��� f%� C�$���B�+\D�wSB�����\~<sv��[q�SQ�c�E��^���^7¾E�,�{�ݡ4}�BF�6r�Ǵ�(����=j����.�<�aoٌwBS�)ƶR������8Qd����J�����SIH��{-�ߦ����"i���o�:߳����,!F�T�<�E�ɨU���`|��Z�n V'g�Zpx����7��r0�.Z�u�DR_�S���Qd��kʯ�}�H����4�r%��dL˓�܂j�ͥ�RomHG��gli�C�xd�����ލ��9��H��?J�'������KQ���kw{5�ᴫu�ҮÃ��}Y4[v8q�\�#`{���ڋ�6�)�K���LjG�Q}�a���8ڄ �DRed���ӷpx%��~:��˚{�������^<;�&֭���+�ł�g�Lȟ��1r�sᙝ+^��`P��������̈́�������ֿb⤍^�rl�>�zz�P+��!%����댂�Hv��h<z��Կ���.l��jo�RQ'�#[���N����}]M�*z��}�͖M��Q�N�d�K�P8�zO�H�/��9�xw��*H��XS7`B��4���fw�Ί�r�;w�Z����9J:�L�3�^�I�׷�/�U�]V� ���#�o�^����$��<R��}�:��.����j��&>aA`c�Ę�w���$:�_�l�_F�֝�m�YU�=��we����*K	�����0G�d�p����H���n�Q���3�r�Tڕ.Mh�d�޿[�2�6��)[�;P����9%���f���y7/��۹���S�8B��X�v��5��)��Uqv���Y�y�pHu;r���辍�q̾xw�>,o��}�b~��O�mE�����}J�"���3�����G�m-W{g��Kml�C��:aef�+��Ɠ&�8�rG��wxϳ���~�A1��uTw��R��i���$v>r�]�m��q��4ݥ*?w�O�=���*B�u�9��d����ͺ�v�_����	���3=�$G�V+7���
�͘��&rD�s��I��(���T�=_��q6��yn��Zm��anۄ��"7��Y�$I�ظ�69$��;�׃���)fA�A&�MtƔ��e�/��+.>��-!�~�Z���Q������]y�E������lX;r��6���H��Z��۪�J�5H�V�u�<
�b��5���abi�zB�R��ԉc�����G�ŕ���6�Ϡ���x�U+r�(Zq�;5��e��-���%R�&�~�jF�\����W)Lp�Yh@����=�gb���/�<���ȼ�}����h�p˂UbU
�97� ���D�"����FΉ=�%���⇋�ڢEɟ�	���O"�Ԧ5�Fe�Y�;��޻É�W��T̆-ǩ�Nd��)m�ެꁞ�+`E���ήc5˪V"cKs�V�����-/�bj3�Գ_����=m�X+��lw$�F,���>1Ŀ��F*��r���{V�VS�����sbk[A�u������As����e:w:l�R���ɱn�҇�"�mr�f��K�M��ݒ�ק��1�D��@�߂M�ӊ�X���2li㛿����.�_��M3_��P�?=#$�P�4~��q�	x����K����T����P^l�2�SN[�6�l�ʶm�pKe��zn�-V `����k�j���wn����Bfa���ھ}�e<�ժ��]�f8�m��B��̂G����z𗫆�$����|Ǣж %�w��o�N?��v�RSҜ&W��,���l�sV�>��iq���8TߙO��G��w#�p����f����)s�zG�� �)%���r�����<��������v7�
�_���{������#3j@a���p��e����"��ၓ/<�}���t�0���~j�^~��l��YJ�6�A�]4��X��V!��V����2�	e{�ᰟJmX�4e��"x�q����ۻ��awZѬNB�������p ;��b�*�#��[1��s�8��5J��D�;�n܏��2)|'�N�L�ץ��bmɡ�B�(�w�v	��	��R#pV��;��Y�v�hwzE�Re������BZA�6�\CF�����?7ʮƷ]Q��gM��}�0�|K�<YR1�;�4���!����O	��&���\���1Ս��S�{'�4'�.��J�Pޠ�c�]�E�Q(�HN2��؟�^C��|��f.7	P#A���Z��N'V��8��Z�(-�NZN�W��u�Шw�ni츑W+��y�I��F��[�+g��L�J��X�ǻ�������]�6,�����-1���Bw������%@�����<"�����t"�ۆ[Q|/�[�^x���/�,�Z�V�|4�I��b��Qnv5;a�?�/�x���=���VN���s��5�W��I��峬8�F=w�F^��yG�3=Q��?�Y_K����p�D�'< ��l�bۗ,�Llmz(�����O����r���ڳT3e���9m�R�}3������*��7��v�:��#SH�o��5I6$vj���Y�� ���AZ���qqH�9��D!(^9�a0����&��I���i�MM���%Z�後S��
g��NfL�1�ͻ�vB���48
3��T?���+�T���a��F)\_���F�J7汖s#���y\Il��X�|����8�w�-`�θX��n?YIU�,��'�F��K2��Z��'���h}L߁�g 
�w��-����Z,������dw�b�p�9'QS����7	c[;c剤��'��6ۓ��ȼLf�j�`RUB�b'�T��w�{��� W�^S4z�|=jZ�xX<5��K)W|6��4�4������ć����>�V����Gpx��d	������6ĩ+�\���s�������H��6�a�*Kī��((��R^d�r��4��y��Te��Sس�eR�F�im�OR|� �J��(�<��|u�z���ь'�FH*��M71q�:%�`����n���և_zj �:Up\�3T��Q�[����o�!A5�}�8��H�Ab�-#MzC*t��F6��Ӹ��U@d�ku�&&~ �����U\��i���!�Kv���j��=�38F@s�O�&�w�-��8_ǩJ����RE��@��ŷ��sN ��X�=�1C���A�l�E��2kmH|��Зz1���x%�+�� ǗϘ�� �`����~!�G�}�y-㍫.����$7��,%M�O�� ����`
�5�(eY+z,��v짟��ޭy{�7�~������_eh��0՟�w8?��$s�E"J7���x�_���	�r�����+fC4�\io�_�F�>�A�a�F��<��%�XMbUœ1��bp�� ]�������U}it��[���TW�bp ���׫ĭ�3s^�}N���+Zk(�2����F�Zu&�����|`�ǃ���m���Y1��Uc��$��·(�?�+Y{�Օ��N�+n�U �S�u���p��0�:����#54z���˽G�`�zbA=F���q�~x�&�H�),h��m�&��m{��rXw��9�q�;���E�8�0r��NU#��Z.�="�X��@�3�ȞC�u&���F�ڐ-��tu#�:G��w��:���)#�5SX~R��U���T0A�ѕ�)�����q<�N��������|���~��#�!{�f�������P���IĝZ��J�C����򲸿��fL���պ��T�=�cG�������r�g�О���/9�M��ຨ)�8����8����I6����������e�X�؆��L��A��&|I�;�#�$?���-�&��MQ[��t{�(e�vi���ET���9��A��wL�97纟�X�&�.�񮫜ze�msD3����Q��-�*�G@��J�s�4�������J|��qХ=)Q�c�Mo��I��@J�U�9�IL�*�@P.��A��Y"�ȥ�q����l˙����[*Y����z;��}��{1��'ɑhؙ�C�7�y�j���[�@R���]�)�e��Sf�=r���o��� ��e|r�c�"����]5&��� G��O�	��[C(�d�?�G��*��E
P]��>��)0?��j+��=���g�Ș>x�
Y��&��j\2� ���T�f;5��� '�����Ě��o=r:�:�(l�.�WQ��@l=`���i�%6;�Sj�	MZ9���^�?+����&����+�uFhV�r����=}���nX�/���֜9o�62�y�O�'�6��N��P�]�&�ӂ��wk����A�n��w"�dg�6˿�� a}îs����+j�<]�(���\<��}⼢.�<�o�����|�&d�ԧ:l-}��_��Ճ��x�H�Ë�`��&���V"�.�L�Z��@H��f��kM±�a�$\�<{찦��G��� �9��|������J�$m�8�t��{p�(G`5*��Ѳ��v��,��p_@�+����@�ȌPe��h�G.5V���ׇ�� M���0�d&%��Z7�[��R{�ɇ����&~_����H�VQX�Ã�o2�%�Pj�Gn�*���d��+P>���X8�ͳ��(��g��;��2�P��yW��f����B���+�2��%�1�X�D�I��]D~ߥj_�x�؏��>�s��� ~�Hv}���,f������B�8�>�؝+ {�Nؿ_�{Ҟm��g_�N+Eb=/��i�I@o�&^{�WE�.����d��t�@�����u��$xc�C�*��A�������6�~u~�����p�_��dr]C��!�l���g���"ۤ���s�L7���	��L��?��۴�3��'񧣶�ה1�R�����M\�tr�X�������L�t�-��=�rvt���SSPn��<n
��#D��p�*(d>	�{��6�iK� T`����r�>��C#�����M��������ZK�1�ž�"�� m��i�H��u�{�}/�A8w*��ixl3����5t�L�'Ja��O���܍��	3�t �3����PSM�o�>�_U�{����a�	qA@��]X���V�1�T��c�3�W�B��q�u�"�>���	�׹F镗UU�a��69e��;� +�
��C�H��/�f�ݲ�lv����{x��7N!屩[�l-��W��JH�cS�:j��W_�%'��E9�')��^p�L�z8�R����7ı8�q�N���w��y�x-#v�M�P��L����;�o"P�:,1� ��������3�����p!Ѷ��Ri����
�Qd�Oȝa��p�}����8�y�bQE��Ƭ���k���p+�,�[W,u��G�����h��7���6��j⟻�=��a�]f�o(gS.ו �#�N�9�z��m���ץB��0%�j�Q�s�����F���,�<�N��Aܑ[�TG1N4B����j+�_׎mC�L��Y���,�q,�����!�KL!��ln�g�<��A���3U�p����+�s��(�R�_
ۧ��F���VMKC�8�!?���}�h?�¼�<�XK��4��!w��T�s�g�H*���A5dD�G=r�L<���l��!�5M�J�p�Z�O�=�!c��m�91�iR�u�{�H��-���'�EjJy�Bn�Ć��aB'6����چ��J?v%���,�	���~��?��e6w������v���BO&�:�����m��ɟ����dP\UD��[k.��nM����G�=\<5te�w�r����}�lzQ"	8��������ۘ�(g�}�.����
�5O���ME��Xkb\�V�����.k���o��Mǜ��� u35D��5�����ۣ��Cy��HJsl��N�	�J�z�8�џfopZt ����^�_"�ݣwL�d��V��٢�}�޵����8+�/�^ܝ��J˃������g��	ym�4�բ�i��#��tg?h��f�B���*kϩ������	�z������JF��5,�|e���="��>_�/g:��eo�g)v,q�H�>���:�x�h���ܴ�f���3�.�H�R�9���5X���<h����gD��s&�(I ������)!��k�^��Y���9)�y�,���0I=�"->ijV���2����eBx�������S��B�Z���W+�X@@�\c˿���[6��)�½�4��r1��6�Λ�E���ď�w;,@�w��p��k1'�I�����ǩp����ǵ!�3@��B��X���b ϛ`�_T�Éy��;��xe��t`�0��Fn�p��xP����p�d�B�
<j�8A��wX�Ӫ4D��^a�E�Ν���P�$������ ����^9�-
\t���iR�(D�<+�_T�f���%�H��fncR�Ŋ+��4���Ƭ:�=<`O�B�<O9��a�Bg�,��g�X�.�;O�=jd;�5����d@��n�d!9EXk��r�3������8n��[��5=���K0����*��´D>���tKY(]�旦����� >A�99��څ�o��ߨ��[(�!���o���߬��.��B<vb#4�_ꃇRC;��U����?[����:��T���:#.�"��ߤZ�H㣅P+��d��ٖ�f�D�͸�������������Q�#L,У�Bz�B���t�\�q?қT�6O����W�r.�nNA;�//--l���������K�*ƙ$Gn@��;-D���G�+_I/�XC}�W����E40`��uy=�7!�Ub�'��Yb�����_BK��ߝ��vr^�+H6k"p�B]��MY�A�Lc�r�1�|6KQ����?1$�!Q���D�찓�]5v�7Hp��ة�����l�;�fqw:���5y�
	�w�[��,�s��O��sBw}d�l��t���{�x��q�t���e�d#sӼ,)��go����n��F������ej��O� �p:g��s'�I:�t���K"�<DQ�"��!��J���4��J\������N�q�'��rֻQ\�m����?�:����:�`5�k1�U����e���\;�S!�S�P:	�4���n0K���ZX�:��U�&�"}��[�;ئ�%<C����s�1{�;��{߉Ž�nl��U7.�s����zk�*���(=�I/�\�\X��T�`@�8���[v��aV*��P3Ť�/9��"/Vfr���['��:MC�@��`�z��v�g�@��=��4���n�u+]�4c���m�qU�a��8]�h���z�bPF����~�GM,W]>Q��/��mgN�̀c*����uђ����V�5)�[�*y���ǒ�H�ZOeWF8�L�~���a���-6Y�ubMs��]
z�z<��F�a�*֠m_q����"�=��BL?�83�]�bƠ�{��|��^AJ ��}�O������k	�ժ�L�!B��	�����3����'�y޸�XP�����e�w�u7+��n�w���% ��b������T���1�&ث%8�9�(�i�	d��|K��L�Ǚ��#75<h�b���%Z�:ЬSf�����_�lH+d#�{�Ej�ԙV��l*<z�M/�q�{
�0�� �TQ��@���)c<%vh9h�P��J�H�l�:���1��L&�9�]<S:8�X]�qF��5�䤙�� ��7$�s���_��~t�%͂O Ʉ�Y(~u^�o���X�p��N=v섡��]�B�r]�F�.$q9�F�Pok\8y�{ȟ�
f�V>/:�Y��?���ǨI)4H�|b�H�XC!��,!ڴ	�7<U��2~�O��M�º��}m��a�`����p��!��;�p����<�Q]8	j�i�pĉ�Xo�mm�$"�Ȁ[��X�:TC.����]M���ͽun2�§�O��P��n.��k(�Y�)�i\��2v� �a_xwC�K�p�q�g@�Od.�|iM3tG�������Nw�0�R}�N��tO�at+5��<���oL�T�6I��f����Pj���Cs����R@b�D��/:]Cy;a��Ǧ��+��N?�u�)G�\�o�K�{ �*�zo��o<�#z��I�G�ٲjv�1~Omt�`�ǩ���)�:&�M�,͑+��g<�%�U *���BF�C����)����+�&�c�-�ƿ�\��|⠊\1��QU�;n�i��"9K��'�����|��5� h� Xy�q�d��6�4 g�L�0A�� v������~GX}0�4���o���"K�â���A4�1G'���G/С}�ʾ�B��B�x�m�h�h�k/m(��%��W!	%�P2gyLj�Wr��#��v��5�b)ه���n:�?~�fpf�bM��F0�#���u���-J�W��Dyj�B,
`�g���7���S	�����P��)Z�E {B�畀��:ɥ�U�g�)28���n֔���y������G�� ��Crp�1B�[6�j�BQ�-�2&P�L�X�Մ�O�>a�T�Q���*)�[���?5U�	0�2���!��g&J��u¾�SNOӫB8��ċ�9P�i�� 1?_Ĥ	X�7!{s��w^��V�@���z��!�GYΣ�� �);�C3��y|	P���ӣ�ۮ�Ņ��c�k�74xV�V�	>OU|��]ch�O���au����Q�P���qe!��ͼݶ����v�7V���:Z���_?��oW1U���!�2]���@~>����(��#��?4��(t&V�m�:[���=P�o��!��
�8tە�`��\��r�>���L�0S�5�s�B2`̘+���A��G��lise�FC�M�fx������Ԯui$5Ż�A�,�9���m�'J�=kO,}J���[�<g�H]�L��e�ӝ t3/��N�P�i�JG�5�A�����>�p�3�\c�t#hU�5�0jc����7��䙇U\�`�����6V)XM���`�9A�(�F
w�=Q�-�ć�"�zԦ���}}��$�[w�,�|;-a���iO.�=1�ě�*u�d�ꔿ�Fh�K��A ��Pn�<��rj�j��	Ԇ�>��o���M�qė�­�]�{�rOb,�SKoo+�@mG�wt�m�&�!7PR�"������ž"�>܋V��Ht>ԹKX7�����3�w�!5<�T&��{�9��u�P=��T�(*�I/>B{��˧6w���a5�[d�/
��  �2�m��n>�?lDu%i��iY�O	�MK3��@���V�]�f�/�C��"H��pI����oW��ę��'h�?f�[i��?��:Rg�g�=+ԧ���|�E��S�zNr�N�5%  1��m�ι�-��t!��|6ů�Xy���鴘	��i�S|�U� 
3�;��;�,]I�1�%.��V�P} ��e����}�Q8�(�� ���	.��9�G�ԥo��Λ�7.,���Z�`�8h�謳�B1�'�1_��vX����`��K��z�'H���Ѥ�/X���y3�)�<h�dTo��U��V5>o��V�嘉���K��(v�m|2ʘ_�i�m�;ۙ�װM�|s�
�,\���*���6�`�����f��Pmt�w�
� �_	��ܞ���V�4y��hBe&J����vM��<��E
y�͏������/fn���?�}��(3�m�,���]��ZF�m��Xښ��<�z�٥������9/��a�}p.I��槐�l�)>Ⰴ{�S\�v6}vG��0_!��״�6��O])�M�#�;�M����!߿!�(������*.5%~_��Ecy:�p��G���\�Bvp�ƚl:�I��R���ܨ[p�T��!�T��x�[��kҙ�q�T���^o�{����i9�O�������dpJ�1��H�f�[b*[`�mB8X��͉\t�U�\�`��^񰒨�$����R�_����yJ���f���.��@�ĺ��
��cw��=΂���W)I巸�~@����`�G�S���zb
���ʠn/���Q}�А�)ILz�/P�d��[q�[���.*�8Lr���>\߆S���
�E�?���9r��7��0XYV���H���{�!>�&%�]{d��$$V�z�2�޻{b��/9��w�Z�;g��4�Y!��[y�C��M]i���͆�BW�\M�x�r�kz�6�k��1�=����[��R���t��߃l�ۆ�s���:-n�P���+�2[��6�o�
��(���<U���DN�(�J~.��E]Rܷ8��[� ��@��a�	���%fC�jj���>�j+�6e0�n��>G�W�ICǄiz�/3v�F��K��yT̖x4q����jS��8v��xo�y�(W�ps/R�vS=��~U"�6�qon���g���DT�7�������8e/HC9m��D%�����;Hԫ&���{[���7��
��O�Om���B����9�j�%�o�ˠ�^`f�t�L��YmzP��k��\F�ڐ����%��|(<A�mԧ?�S�P/D�C���RU���$;x�GT��}	�"�Z�UA��w�(�G�t���?���DS��� 7]Gz��~U�J�#��P���f�[X,}ؤFL3�B7h=1�Q��h�jf��C���+Q���[��J�ع�������C2!�m'�D{����d��n�*l�ۿ�������y�"*#�����֐�s�}���z|R�{�c-���XA�ŏ��(;!1���_���oN�d7��8L���������1m�."��5G�X7��wL|w㖵�Cp��2k�@(
�''Kv�c?�J���o�G�;�mZrc'�%&!5�HjyL�2�]���{�����8tfvlX�(w����|~�|<�+{�q%�7�(N9ؕ����/�lߨ�#��������'T��X���Ԋ�=v�7�'FcAo�r|gԨEfL/U[�t���}��n�]�AUu\��{��W1�#W�uX.E���0]R.�y�S:��7k�}P�5n��Ԇ}_�m9�Uu�]_'�umC��3&~U0��ŀq���"Iꑐ賚b����R�I����͆v�=��ia��ʧ�L�.y�p��g�޽*�s��!�M��[�a�x(d��XIÝZ�s�'{_���C/�Z)_����F�r?`b;�T8���r�%(�)�sQeEu�i�� 66��ri%�0������_�E����8\q�$K�]�Pw�l�]���W�A�x-���o�*h��3���=JwQ��iP�UQ���VoRW�wa色�8��.��JM������O#��Y�Qo�6��X4��o���Y,��C�%��W��?%C7b)�� �r� YF�0{Zj����~�y���$��tNtR��X/g���Ƭjr�e��:������{z���/�k��{³���@I�^�JA�]��#J��BFl��q��4m����q������[�Inb�-��Nq6ο�V�����Y˘z�y�� ������ӊ��3U�;��w*�nl�Z���i��;�'���!�,�.$f����C-�g�L����bjN��~Z�A�@�p���x���*p%]�Z�9�BE����z6)ȸ��(ޗz�U0]��oZ���fWBg�*��ڛk���pqk�5�אh��FO��q�d�cP�5 �I����;��J�;��)���j=:p�8�!(>�n�^S�%�3�@� �V�f��]l9
��B%'�:2S2V���|�a�\���tkQV��z�Ai��3��1�E .����7L�~�w�?���Mon�6# �C�O����%�+���-�֓i)��D��y��t�0u�H,۽�t0g�<v�VX?s�uI��>�҆��"�Yà0����m��`�̏���z��0"��ʇ3(��]!?ȱ7�2
�2,�$�늚a������9�6��]� /\��zp��lp����)�Fe[s>�2$�~��neJ��8�BѠ~���
w݅+�\���Z�o3���"�X��']C�M�À*4��;�IO��_��W1������m%�;(G�Q��X�_�<���!��^J��>RJ�)?�t�X�k�e���US��2 x�����<r��y�/��\��A�4=��i3a)��F.h��t�g�ez�ks�K��f�P��!�	�Q@�-�	LouL���h�,�z�I�����|�6�%E,fV^�D���Ğ5d�L*�P�1�:�TK�7��|$�W>:Q>i-G�8/�ÈV�BTS�ss��M����M�oZ���,�p�,xz�v���Q���߾`r�4"����Q`W�5�]�/!�c��OZ�K�	Tn�D�C�.���iP2����0y���G�<s}�/��b�B��PŬ�������ɨg����&8eK��3a����v������o�a�"���6&!7c��B���jg��k�}�N�A��AR�i+Z��E�3c6�QI3W�]����[kB��{����0������Ȁ��	�"��>R��C�h�B��
���-�0S��~�
z���wWF�Ȝ"�������F��+��r5d��0FܽJjW�D^؆��{�V,��e���7R�ggy�fH0��ށ�'y��f��?��͇#i疳Y��'���r��i����)�!AA�W�4oуA���������!?A`�!ˋ�Pb�j�&6�ׂ�~���1���6���v�E��9�!J�r�����$
��.Ů�l&}�ڥŰt�%���S�G7������BpFH ��VY��6��e���=@�Ke!��P�YЛ3y�LK��Q��� ��}���J�X�	{ӊ?�ի��lV�ê��W�P� ��L	��8��ۑ�)����y`�c�j1[�=�{��J��+��(����B�Gy~�N"��:,���NQ���t�աr�p|Tl�J���8�b����8C�R̓��Tr�ƥ8���.;����z��պ�G�3���X��[Eu��UHZ�z�Fc�C�~�ճ���{�����H�y۽�yp�OR��Ѧ�H���q�
$����`.y>JKKa&�l�Q|������{0j��YE��r�`�&��ݡ����xT�n=� v&yNI%mRY�3Xz���og2o4��!��V0	�qc�����"�W�:�����a�(��~